magic
tech scmos
timestamp 1492460222
<< metal1 >>
rect -112 1150 -106 1154
rect -66 1142 -50 1146
rect -112 1040 -106 1044
rect -66 1032 -58 1036
rect -112 930 -106 934
rect -46 930 -42 934
rect -66 922 -50 926
rect -2 922 6 926
rect -112 820 -106 824
rect -54 820 -38 824
rect -66 812 -58 816
rect -2 812 6 816
rect 46 812 57 816
rect -112 710 -106 714
rect -46 710 -42 714
rect -66 702 -50 706
rect -2 702 6 706
rect 50 702 57 706
rect -112 600 -106 604
rect -54 600 -38 604
rect -66 592 -58 596
rect -2 592 6 596
rect 50 592 57 596
rect -112 490 -106 494
rect -46 490 -42 494
rect -66 482 -50 486
rect -2 482 6 486
rect 50 482 57 486
rect -112 380 -106 384
rect -54 380 -38 384
rect -66 372 -58 376
rect -2 372 6 376
rect 50 372 57 376
rect -112 270 -106 274
rect -46 270 -42 274
rect -66 262 -50 266
rect -2 262 6 266
rect 50 262 57 266
rect -112 160 -106 164
rect -54 160 -38 164
rect -2 152 6 156
rect 50 152 57 156
rect -52 90 -43 98
rect -112 50 -106 54
rect -46 50 -42 54
rect 50 42 57 46
rect -53 0 -44 8
<< m2contact >>
rect -50 1142 -46 1146
rect -58 1032 -54 1036
rect -50 930 -46 934
rect -50 922 -46 926
rect 6 922 10 926
rect -58 820 -54 824
rect -58 812 -54 816
rect 6 812 10 816
rect -50 710 -46 714
rect -50 702 -46 706
rect 6 702 10 706
rect -58 600 -54 604
rect -58 592 -54 596
rect 6 592 10 596
rect -50 490 -46 494
rect -50 482 -46 486
rect 6 482 10 486
rect -58 380 -54 384
rect -58 372 -54 376
rect 6 372 10 376
rect -50 270 -46 274
rect -50 262 -46 266
rect 6 262 10 266
rect -58 160 -54 164
rect 6 152 10 156
rect -50 50 -46 54
<< metal2 >>
rect -98 50 -94 1208
rect -82 59 -78 1208
rect -74 1145 -70 1152
rect -74 1035 -70 1042
rect -74 925 -70 932
rect -66 915 -62 926
rect -58 824 -54 1032
rect -50 934 -46 1142
rect -74 815 -70 822
rect -66 805 -62 816
rect -74 705 -70 712
rect -66 695 -62 706
rect -58 604 -54 812
rect -50 714 -46 922
rect -74 595 -70 602
rect -66 585 -62 596
rect -74 485 -70 492
rect -66 475 -62 486
rect -58 384 -54 592
rect -50 494 -46 702
rect -74 375 -70 382
rect -66 365 -62 376
rect -74 265 -70 272
rect -66 255 -62 266
rect -58 164 -54 372
rect -50 274 -46 482
rect -74 155 -70 162
rect -66 145 -62 156
rect -50 54 -46 262
rect -74 45 -70 52
rect -34 50 -30 989
rect -18 59 -14 989
rect -10 915 -6 932
rect -10 805 -6 822
rect 6 820 10 922
rect -10 695 -6 712
rect 6 710 10 812
rect -10 585 -6 602
rect 6 600 10 702
rect -10 475 -6 492
rect 6 490 10 592
rect -10 365 -6 382
rect 6 380 10 482
rect -10 255 -6 272
rect 6 270 10 372
rect -10 145 -6 162
rect 6 160 10 262
rect -66 35 -62 46
rect -10 35 -6 52
rect 6 50 10 152
rect 14 50 18 880
rect 30 59 34 880
rect 38 816 42 822
rect 38 706 42 712
rect 38 596 42 602
rect 38 486 42 492
rect 38 376 42 382
rect 38 266 42 272
rect 38 156 42 162
rect 38 46 42 52
<< m3contact >>
rect -74 1141 -70 1145
rect -74 1031 -70 1035
rect -74 921 -70 925
rect -66 911 -62 915
rect -74 811 -70 815
rect -66 801 -62 805
rect -74 701 -70 705
rect -66 691 -62 695
rect -74 591 -70 595
rect -66 581 -62 585
rect -74 481 -70 485
rect -66 471 -62 475
rect -74 371 -70 375
rect -66 361 -62 365
rect -74 261 -70 265
rect -66 251 -62 255
rect -74 151 -70 155
rect -66 141 -62 145
rect -10 911 -6 915
rect -10 801 -6 805
rect 6 812 10 816
rect -10 691 -6 695
rect 6 702 10 706
rect -10 581 -6 585
rect 6 592 10 596
rect -10 471 -6 475
rect 6 482 10 486
rect -10 361 -6 365
rect 6 372 10 376
rect -10 251 -6 255
rect 6 262 10 266
rect -10 141 -6 145
rect 6 152 10 156
rect -74 41 -70 45
rect -66 31 -62 35
rect 38 812 42 816
rect 38 702 42 706
rect 38 592 42 596
rect 38 482 42 486
rect 38 372 42 376
rect 38 262 42 266
rect 38 152 42 156
rect -2 42 2 46
rect 38 42 42 46
rect -10 31 -6 35
<< metal3 >>
rect -112 1145 -69 1146
rect -112 1141 -74 1145
rect -70 1141 -69 1145
rect -112 1140 -69 1141
rect -112 1035 -69 1036
rect -112 1031 -74 1035
rect -70 1031 -69 1035
rect -112 1030 -69 1031
rect -112 925 -69 926
rect -112 921 -74 925
rect -70 921 -69 925
rect -112 920 -69 921
rect -67 915 -5 916
rect -67 911 -66 915
rect -62 911 -10 915
rect -6 911 -5 915
rect -67 910 -5 911
rect 5 816 43 817
rect -112 815 -69 816
rect -112 811 -74 815
rect -70 811 -69 815
rect 5 812 6 816
rect 10 812 38 816
rect 42 812 43 816
rect 5 811 43 812
rect -112 810 -69 811
rect -67 805 -5 806
rect -67 801 -66 805
rect -62 801 -10 805
rect -6 801 -5 805
rect -67 800 -5 801
rect 5 706 43 707
rect -112 705 -69 706
rect -112 701 -74 705
rect -70 701 -69 705
rect 5 702 6 706
rect 10 702 38 706
rect 42 702 43 706
rect 5 701 43 702
rect -112 700 -69 701
rect -67 695 -5 696
rect -67 691 -66 695
rect -62 691 -10 695
rect -6 691 -5 695
rect -67 690 -5 691
rect 5 596 43 597
rect -112 595 -69 596
rect -112 591 -74 595
rect -70 591 -69 595
rect 5 592 6 596
rect 10 592 38 596
rect 42 592 43 596
rect 5 591 43 592
rect -112 590 -69 591
rect -67 585 -5 586
rect -67 581 -66 585
rect -62 581 -10 585
rect -6 581 -5 585
rect -67 580 -5 581
rect 5 486 43 487
rect -112 485 -69 486
rect -112 481 -74 485
rect -70 481 -69 485
rect 5 482 6 486
rect 10 482 38 486
rect 42 482 43 486
rect 5 481 43 482
rect -112 480 -69 481
rect -67 475 -5 476
rect -67 471 -66 475
rect -62 471 -10 475
rect -6 471 -5 475
rect -67 470 -5 471
rect 5 376 43 377
rect -112 375 -69 376
rect -112 371 -74 375
rect -70 371 -69 375
rect 5 372 6 376
rect 10 372 38 376
rect 42 372 43 376
rect 5 371 43 372
rect -112 370 -69 371
rect -67 365 -5 366
rect -67 361 -66 365
rect -62 361 -10 365
rect -6 361 -5 365
rect -67 360 -5 361
rect 5 266 43 267
rect -112 265 -69 266
rect -112 261 -74 265
rect -70 261 -69 265
rect 5 262 6 266
rect 10 262 38 266
rect 42 262 43 266
rect 5 261 43 262
rect -112 260 -69 261
rect -67 255 -5 256
rect -67 251 -66 255
rect -62 251 -10 255
rect -6 251 -5 255
rect -67 250 -5 251
rect 5 156 43 157
rect -112 155 -69 156
rect -112 151 -74 155
rect -70 151 -69 155
rect 5 152 6 156
rect 10 152 38 156
rect 42 152 43 156
rect 5 151 43 152
rect -112 150 -69 151
rect -67 145 -5 146
rect -67 141 -66 145
rect -62 141 -10 145
rect -6 141 -5 145
rect -67 140 -5 141
rect -3 46 43 47
rect -112 45 -69 46
rect -112 41 -74 45
rect -70 41 -69 45
rect -3 42 -2 46
rect 2 42 38 46
rect 42 42 43 46
rect -3 41 43 42
rect -112 40 -69 41
rect -67 35 -5 36
rect -67 31 -66 35
rect -62 31 -10 35
rect -6 31 -5 35
rect -67 30 -5 31
use mux2_dp_1x  mux2_dp_1x_6
timestamp 1484435125
transform 1 0 -106 0 1 1104
box -6 -4 50 96
use mux2_dp_1x  mux2_dp_1x_5
timestamp 1484435125
transform 1 0 -106 0 1 994
box -6 -4 50 96
use mux2_dp_1x  mux2_dp_1x_4
timestamp 1484435125
transform 1 0 -106 0 1 884
box -6 -4 50 96
use mux2_dp_1x  mux2_dp_1x_3
timestamp 1484435125
transform 1 0 -42 0 1 884
box -6 -4 50 96
use mux2_dp_1x  mux2_dp_1x_2
array 1 1 56 1 8 110
timestamp 1484435125
transform 1 0 -106 0 1 4
box -6 -4 50 96
use mux2_dp_1x  mux2_dp_1x_1
array 1 1 56 1 8 110
timestamp 1484435125
transform 1 0 -42 0 1 4
box -6 -4 50 96
use mux2_dp_1x  mux2_dp_1x_0
array 1 1 56 1 8 110
timestamp 1484435125
transform 1 0 6 0 1 4
box -6 -4 50 96
<< labels >>
rlabel metal2 32 878 32 878 1 s0
rlabel metal2 16 878 16 878 1 s0b
rlabel metal2 -16 987 -16 987 1 s1
rlabel metal2 -32 987 -32 987 1 s1b
rlabel metal2 -80 1206 -80 1206 5 s2
rlabel metal2 -96 1206 -96 1206 5 s2b
rlabel metal1 55 44 55 44 1 y0
rlabel metal1 55 154 55 154 1 y1
rlabel metal1 55 264 55 264 1 y2
rlabel metal1 55 374 55 374 1 y3
rlabel metal1 55 484 55 484 1 y4
rlabel metal1 55 594 55 594 1 y5
rlabel metal1 55 704 55 704 1 y6
rlabel metal1 55 814 55 814 7 y7
rlabel metal3 -110 1143 -110 1143 3 z10
rlabel metal1 -111 1152 -111 1152 3 z14
rlabel metal1 -110 1042 -110 1042 3 z13
rlabel metal1 -110 932 -110 932 3 z12
rlabel metal1 -110 822 -110 822 3 z11
rlabel metal1 -110 712 -110 712 3 z10
rlabel metal1 -110 602 -110 602 3 z9
rlabel metal1 -111 492 -111 492 3 z8
rlabel metal1 -111 382 -111 382 3 z7
rlabel metal1 -110 272 -110 272 3 z6
rlabel metal1 -110 162 -110 162 3 z5
rlabel metal1 -110 52 -110 52 3 z4
rlabel metal3 -110 43 -110 43 3 z0
rlabel metal3 -110 153 -110 153 3 z1
rlabel metal3 -110 263 -110 263 3 z2
rlabel metal3 -110 373 -110 373 3 z3
rlabel metal3 -111 483 -111 483 3 z4
rlabel metal3 -110 593 -110 593 3 z5
rlabel metal3 -110 703 -110 703 3 z6
rlabel metal3 -110 813 -110 813 3 z7
rlabel metal3 -110 923 -110 923 3 z8
rlabel metal3 -109 1033 -109 1033 3 z9
<< end >>
