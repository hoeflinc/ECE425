magic
tech scmos
timestamp 1490727808
<< m2contact >>
rect -7 -2 7 2
<< end >>
