magic
tech scmos
timestamp 1493147875
<< m2contact >>
rect -7 -2 7 2
<< end >>
