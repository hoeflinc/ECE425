magic
tech scmos
timestamp 1492457336
<< nwell >>
rect -6 40 74 96
<< ntransistor >>
rect 7 8 9 14
rect 15 8 17 14
rect 20 8 22 14
rect 28 8 30 14
rect 33 8 35 14
rect 41 8 43 14
rect 61 8 63 22
<< ptransistor >>
rect 7 73 9 82
rect 15 73 17 82
rect 20 73 22 82
rect 28 73 30 82
rect 33 73 35 82
rect 41 73 43 82
rect 61 62 63 82
<< ndiffusion >>
rect 2 13 7 14
rect 6 9 7 13
rect 2 8 7 9
rect 9 8 10 14
rect 14 8 15 14
rect 17 8 20 14
rect 22 8 23 14
rect 27 8 28 14
rect 30 8 33 14
rect 35 8 36 14
rect 40 8 41 14
rect 43 8 44 14
rect 60 8 61 22
rect 63 8 64 22
<< pdiffusion >>
rect 6 73 7 82
rect 9 73 10 82
rect 14 73 15 82
rect 17 73 20 82
rect 22 73 23 82
rect 27 73 28 82
rect 30 73 33 82
rect 35 73 36 82
rect 40 73 41 82
rect 43 73 44 82
rect 60 62 61 82
rect 63 62 64 82
<< ndcontact >>
rect 2 9 6 13
rect 10 8 14 14
rect 23 8 27 14
rect 36 8 40 14
rect 44 8 48 14
rect 56 8 60 22
rect 64 8 68 22
<< pdcontact >>
rect 2 73 6 82
rect 10 73 14 82
rect 23 73 27 82
rect 36 73 40 82
rect 44 73 48 82
rect 56 62 60 82
rect 64 62 68 82
<< psubstratepcontact >>
rect 0 -2 4 2
rect 8 -2 12 2
rect 16 -2 20 2
rect 24 -2 28 2
rect 32 -2 36 2
rect 40 -2 44 2
rect 48 -2 52 2
rect 56 -2 60 2
rect 64 -2 68 2
<< nsubstratencontact >>
rect 0 88 4 92
rect 8 88 12 92
rect 16 88 20 92
rect 24 88 28 92
rect 32 88 36 92
rect 40 88 44 92
rect 48 88 52 92
rect 56 88 60 92
rect 64 88 68 92
<< polysilicon >>
rect 7 82 9 84
rect 15 82 17 84
rect 20 82 22 84
rect 28 82 30 84
rect 33 82 35 84
rect 41 82 43 84
rect 61 82 63 84
rect 7 72 9 73
rect 15 72 17 73
rect 7 70 17 72
rect 20 72 22 73
rect 20 70 23 72
rect 7 42 9 70
rect 17 46 18 49
rect 7 38 8 42
rect 7 17 9 38
rect 16 28 18 46
rect 21 41 23 70
rect 28 50 30 73
rect 33 58 35 73
rect 41 72 43 73
rect 41 70 46 72
rect 33 57 41 58
rect 33 56 35 57
rect 21 39 27 41
rect 25 36 27 39
rect 16 26 22 28
rect 7 15 17 17
rect 7 14 9 15
rect 15 14 17 15
rect 20 14 22 26
rect 25 17 27 32
rect 39 28 41 57
rect 33 26 41 28
rect 44 36 46 70
rect 61 43 63 62
rect 44 32 45 36
rect 25 15 30 17
rect 28 14 30 15
rect 33 14 35 26
rect 44 17 46 32
rect 61 22 63 39
rect 41 15 46 17
rect 41 14 43 15
rect 7 6 9 8
rect 15 6 17 8
rect 20 6 22 8
rect 28 6 30 8
rect 33 6 35 8
rect 41 6 43 8
rect 61 6 63 8
<< polycontact >>
rect 13 46 17 50
rect 8 38 12 42
rect 35 53 39 57
rect 27 46 31 50
rect 25 32 29 36
rect 59 39 63 43
rect 45 32 49 36
<< metal1 >>
rect -2 92 70 94
rect -2 88 0 92
rect 4 88 8 92
rect 12 88 16 92
rect 20 88 24 92
rect 28 88 32 92
rect 36 88 40 92
rect 44 88 48 92
rect 52 88 56 92
rect 60 88 64 92
rect 68 88 70 92
rect -2 86 70 88
rect 10 82 14 86
rect 36 82 40 86
rect 56 82 60 86
rect 4 53 35 57
rect 17 46 27 50
rect 31 46 48 50
rect 28 39 59 43
rect 29 32 40 36
rect 44 32 45 36
rect 4 13 6 14
rect 2 8 6 9
rect 10 4 14 8
rect 36 4 40 8
rect 56 4 60 8
rect -2 2 70 4
rect -2 -2 0 2
rect 4 -2 8 2
rect 12 -2 16 2
rect 20 -2 24 2
rect 28 -2 32 2
rect 36 -2 40 2
rect 44 -2 48 2
rect 52 -2 56 2
rect 60 -2 64 2
rect 68 -2 70 2
rect -2 -4 70 -2
<< m2contact >>
rect 0 73 2 77
rect 2 73 4 77
rect 24 73 27 77
rect 27 73 28 77
rect 48 73 52 77
rect 64 62 68 66
rect 0 53 4 57
rect 48 46 52 50
rect 8 38 12 42
rect 24 39 28 43
rect 40 32 44 36
rect 0 13 4 14
rect 0 10 2 13
rect 2 10 4 13
rect 24 10 27 14
rect 27 10 28 14
rect 48 10 52 14
rect 64 18 68 22
<< metal2 >>
rect 0 57 4 73
rect 0 14 4 53
rect 24 43 28 73
rect 24 14 28 39
rect 48 50 52 73
rect 48 14 52 46
rect 64 22 68 62
<< labels >>
rlabel metal2 66 34 66 34 1 y
rlabel m2contact 42 34 42 34 1 b
rlabel m2contact 10 40 10 40 1 a
rlabel metal1 -1 90 -1 90 3 Vdd!
rlabel metal1 -1 0 -1 0 2 Gnd!
rlabel m2contact 26 41 26 41 1 yb
<< end >>
