magic
tech scmos
timestamp 1488310061
<< m2contact >>
rect -7 -2 7 2
<< end >>
