magic
tech scmos
timestamp 1493147875
<< m2contact >>
rect -2 -2 2 2
<< end >>
