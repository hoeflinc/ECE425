magic
tech scmos
timestamp 1493692910
<< metal2 >>
rect 487 2552 491 2556
rect 241 1344 245 1845
rect 904 1541 908 1815
rect 924 1719 928 2512
rect 934 1749 938 2530
rect 944 1789 948 2521
rect 1006 2494 1010 2539
rect 1030 2497 1034 2548
rect 1062 2497 1066 2557
rect 1095 2494 1099 2566
rect 1134 2497 1138 2575
rect 1166 2497 1170 2584
rect 250 1380 254 1537
rect 265 1343 269 1523
rect 305 1344 309 1376
rect 942 1354 946 1685
rect 950 1344 954 1645
rect 958 1527 962 1595
rect 966 1424 970 1575
rect 1135 1460 1138 1518
rect 1167 1470 1170 1519
rect 1199 1480 1202 1519
rect 1231 1490 1234 1517
rect 1295 1500 1298 1518
rect 1335 1510 1338 1519
rect 1321 1344 1325 1456
rect 1353 1342 1357 1466
rect 1529 1340 1533 1476
rect 1681 1344 1685 1486
rect 1713 1344 1717 1496
rect 1769 1344 1773 1506
rect 1937 1343 1941 1516
rect 1391 1067 1395 1124
rect 2077 1036 2081 1064
rect 2640 1015 2644 1032
<< m3contact >>
rect 471 2584 475 2588
rect 1166 2584 1170 2588
rect 463 2575 467 2579
rect 1134 2575 1138 2579
rect 455 2566 459 2570
rect 1095 2566 1099 2570
rect 447 2557 451 2561
rect 1062 2557 1066 2561
rect 439 2548 443 2552
rect 1030 2548 1034 2552
rect 431 2539 435 2543
rect 1006 2539 1010 2543
rect 487 2530 491 2534
rect 934 2530 938 2534
rect 671 2521 675 2525
rect 303 2512 307 2516
rect 924 2512 928 2516
rect 241 1845 245 1849
rect 904 1815 908 1819
rect 944 2521 948 2525
rect 944 1785 948 1789
rect 934 1745 938 1749
rect 924 1715 928 1719
rect 250 1537 254 1541
rect 904 1537 908 1541
rect 942 1685 946 1689
rect 250 1376 254 1380
rect 265 1523 269 1527
rect 518 1410 522 1414
rect 526 1400 530 1404
rect 540 1390 544 1394
rect 548 1380 552 1384
rect 305 1376 309 1380
rect 556 1370 560 1374
rect 672 1360 676 1364
rect 942 1350 946 1354
rect 950 1645 954 1649
rect 958 1595 962 1599
rect 958 1523 962 1527
rect 966 1575 970 1579
rect 1366 1516 1370 1520
rect 1937 1516 1941 1520
rect 1335 1506 1339 1510
rect 1769 1506 1773 1510
rect 1295 1496 1299 1500
rect 1713 1496 1717 1500
rect 1231 1486 1235 1490
rect 1681 1486 1685 1490
rect 1199 1476 1203 1480
rect 1529 1476 1533 1480
rect 1167 1466 1171 1470
rect 1353 1466 1357 1470
rect 1135 1456 1139 1460
rect 1321 1456 1325 1460
rect 966 1420 970 1424
rect 950 1340 954 1344
rect 1391 1124 1395 1128
rect 2592 1124 2596 1128
rect 1409 1064 1413 1068
rect 2077 1064 2081 1068
rect 2077 1032 2081 1036
rect 2640 1032 2644 1036
<< metal3 >>
rect 470 2588 1171 2589
rect 470 2584 471 2588
rect 475 2584 1166 2588
rect 1170 2584 1171 2588
rect 470 2583 1171 2584
rect 462 2579 1139 2580
rect 462 2575 463 2579
rect 467 2575 1134 2579
rect 1138 2575 1139 2579
rect 462 2574 1139 2575
rect 454 2570 1100 2571
rect 454 2566 455 2570
rect 459 2566 1095 2570
rect 1099 2566 1100 2570
rect 454 2565 1100 2566
rect 446 2561 1067 2562
rect 446 2557 447 2561
rect 451 2557 1062 2561
rect 1066 2557 1067 2561
rect 446 2556 1067 2557
rect 438 2552 1035 2553
rect 438 2548 439 2552
rect 443 2548 1030 2552
rect 1034 2548 1035 2552
rect 438 2547 1035 2548
rect 430 2543 1011 2544
rect 430 2539 431 2543
rect 435 2539 1006 2543
rect 1010 2539 1011 2543
rect 430 2538 1011 2539
rect 486 2534 939 2535
rect 486 2530 487 2534
rect 491 2530 934 2534
rect 938 2530 939 2534
rect 486 2529 939 2530
rect 670 2525 949 2526
rect 670 2521 671 2525
rect 675 2521 944 2525
rect 948 2521 949 2525
rect 670 2520 949 2521
rect 302 2516 929 2517
rect 302 2512 303 2516
rect 307 2512 924 2516
rect 928 2512 929 2516
rect 302 2511 929 2512
rect 240 1849 965 1850
rect 240 1845 241 1849
rect 245 1845 965 1849
rect 240 1844 965 1845
rect 903 1819 965 1820
rect 903 1815 904 1819
rect 908 1815 965 1819
rect 903 1814 965 1815
rect 943 1789 965 1790
rect 943 1785 944 1789
rect 948 1785 965 1789
rect 943 1784 965 1785
rect 933 1749 966 1750
rect 933 1745 934 1749
rect 938 1745 966 1749
rect 933 1744 966 1745
rect 923 1719 965 1720
rect 923 1715 924 1719
rect 928 1715 965 1719
rect 923 1714 965 1715
rect 941 1689 965 1690
rect 941 1685 942 1689
rect 946 1685 965 1689
rect 941 1684 965 1685
rect 949 1649 965 1650
rect 949 1645 950 1649
rect 954 1645 965 1649
rect 949 1644 965 1645
rect 957 1599 965 1600
rect 957 1595 958 1599
rect 962 1595 965 1599
rect 957 1594 965 1595
rect 965 1579 971 1580
rect 965 1575 966 1579
rect 970 1575 971 1579
rect 965 1574 971 1575
rect 249 1541 909 1542
rect 249 1537 250 1541
rect 254 1537 904 1541
rect 908 1537 909 1541
rect 249 1536 909 1537
rect 264 1527 963 1528
rect 264 1523 265 1527
rect 269 1523 958 1527
rect 962 1523 963 1527
rect 264 1522 963 1523
rect 1365 1520 1942 1521
rect 1365 1516 1366 1520
rect 1370 1516 1937 1520
rect 1941 1516 1942 1520
rect 1365 1515 1942 1516
rect 1334 1510 1774 1511
rect 1334 1506 1335 1510
rect 1339 1506 1769 1510
rect 1773 1506 1774 1510
rect 1334 1505 1774 1506
rect 1294 1500 1718 1501
rect 1294 1496 1295 1500
rect 1299 1496 1713 1500
rect 1717 1496 1718 1500
rect 1294 1495 1718 1496
rect 1230 1490 1686 1491
rect 1230 1486 1231 1490
rect 1235 1486 1681 1490
rect 1685 1486 1686 1490
rect 1230 1485 1686 1486
rect 1198 1480 1534 1481
rect 1198 1476 1199 1480
rect 1203 1476 1529 1480
rect 1533 1476 1534 1480
rect 1198 1475 1534 1476
rect 1166 1470 1358 1471
rect 1166 1466 1167 1470
rect 1171 1466 1353 1470
rect 1357 1466 1358 1470
rect 1166 1465 1358 1466
rect 1134 1460 1326 1461
rect 1134 1456 1135 1460
rect 1139 1456 1321 1460
rect 1325 1456 1326 1460
rect 1134 1455 1326 1456
rect 507 1424 971 1425
rect 507 1420 966 1424
rect 970 1420 971 1424
rect 507 1419 971 1420
rect 249 1380 310 1381
rect 249 1376 250 1380
rect 254 1376 305 1380
rect 309 1376 310 1380
rect 249 1375 310 1376
rect 708 1354 947 1355
rect 708 1350 942 1354
rect 946 1350 947 1354
rect 708 1349 947 1350
rect 712 1344 955 1345
rect 712 1340 950 1344
rect 954 1340 955 1344
rect 712 1339 955 1340
rect 1390 1128 2597 1129
rect 1390 1124 1391 1128
rect 1395 1124 2592 1128
rect 2596 1124 2597 1128
rect 1390 1123 2597 1124
rect 1408 1068 2082 1069
rect 1408 1064 1409 1068
rect 1413 1064 2077 1068
rect 2081 1064 2082 1068
rect 1408 1063 2082 1064
rect 2076 1036 2645 1037
rect 2076 1032 2077 1036
rect 2081 1032 2640 1036
rect 2644 1032 2645 1036
rect 2076 1031 2645 1032
use mips_fsm  mips_fsm_0
timestamp 1493147875
transform 1 0 965 0 1 1517
box 0 0 584 980
use datapath_new  datapath_new_0
timestamp 1493661823
transform 1 0 -279 0 1 32
box 279 -32 3123 2811
<< labels >>
rlabel m3contact 674 1362 674 1362 1 funct_0_
rlabel m3contact 558 1372 558 1372 1 funct_1_
rlabel m3contact 550 1382 550 1382 1 funct_2_
rlabel m3contact 542 1392 542 1392 1 funct_3_
rlabel m3contact 528 1402 528 1402 1 funct_4_
<< end >>
