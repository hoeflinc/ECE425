magic
tech scmos
timestamp 1492976468
<< metal2 >>
rect -33 1621 -27 1622
rect -33 1617 -32 1621
rect -28 1617 -27 1621
rect -33 1616 -27 1617
rect -41 1602 -35 1603
rect -41 1598 -40 1602
rect -36 1598 -35 1602
rect -41 1597 -35 1598
rect -243 1278 -179 1343
rect -123 1308 -119 1312
rect -40 1308 -36 1597
rect -32 1308 -28 1616
rect -25 1572 -19 1573
rect -25 1568 -24 1572
rect -20 1568 -19 1572
rect -25 1567 -19 1568
rect -24 1308 -20 1567
rect 0 1308 4 1312
rect 56 1308 60 1312
rect 184 1308 188 1312
rect 192 1308 196 1312
rect 200 1308 204 1312
rect 208 1308 212 1312
rect 216 1308 220 1312
rect 224 1308 228 1312
rect 240 1308 244 1312
rect 424 1308 428 1312
rect 584 1308 588 1312
rect 696 1308 700 1312
rect 728 1308 732 1312
rect 736 1308 740 1312
rect 744 1308 748 1312
rect 752 1308 756 1312
rect 792 1308 796 1312
rect 960 1308 964 1312
rect 1600 1308 1604 1312
rect 1632 1308 1636 1312
rect 1808 1308 1812 1312
rect 1960 1308 1964 1312
rect 1992 1308 1996 1312
rect 2048 1308 2052 1312
rect 2216 1308 2220 1312
rect 2240 1308 2244 1312
rect 2480 1308 2484 1312
rect 2512 1308 2516 1312
rect 2634 1278 2698 1862
rect 2724 1278 2788 1863
<< m3contact >>
rect -32 1617 -28 1621
rect -40 1598 -36 1602
rect -24 1568 -20 1572
<< metal3 >>
rect -63 1621 -27 1622
rect -63 1617 -32 1621
rect -28 1617 -27 1621
rect -63 1616 -27 1617
rect -63 1602 -35 1603
rect -63 1598 -40 1602
rect -36 1598 -35 1602
rect -63 1597 -35 1598
rect -63 1572 -19 1573
rect -63 1568 -24 1572
rect -20 1568 -19 1572
rect -63 1567 -19 1568
use controller  controller_0
timestamp 1492976468
transform 1 0 0 0 1 1450
box -243 -172 2788 368
use datapath  datapath_0
timestamp 1492976468
transform 1 0 0 0 1 0
box -243 -32 2788 1343
<< end >>
