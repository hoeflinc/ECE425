magic
tech scmos
timestamp 1493745683
<< m2contact >>
rect -7 -2 7 2
<< end >>
