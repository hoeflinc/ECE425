magic
tech scmos
timestamp 1492476009
<< metal1 >>
rect -26 1477 -8 1481
rect -26 1367 -15 1371
rect -26 1257 -22 1261
rect -4 1040 1 1044
rect -11 930 0 934
rect -18 820 0 824
rect -25 710 0 714
rect -4 490 0 494
rect -11 380 0 384
rect -18 270 1 274
rect -25 160 1 164
<< m2contact >>
rect -28 1582 -24 1586
rect -8 1477 -4 1481
rect -15 1367 -11 1371
rect -22 1257 -18 1261
rect -29 1147 -25 1151
rect -1 1150 3 1154
rect -8 1040 -4 1044
rect -47 1030 -43 1034
rect -15 930 -11 934
rect -47 920 -43 924
rect -22 820 -18 824
rect -47 810 -43 814
rect -29 710 -25 714
rect -1 600 3 604
rect -8 490 -4 494
rect -15 380 -11 384
rect -22 270 -18 274
rect -29 160 -25 164
rect -1 50 3 54
<< metal2 >>
rect -28 1519 -24 1582
rect -2 1528 2 1563
rect -29 1145 -25 1147
rect -29 714 -25 1141
rect -22 824 -18 1257
rect -15 934 -11 1367
rect -8 1044 -4 1477
rect -1 1154 3 1515
rect 14 1324 18 1524
rect 14 1252 18 1320
rect 46 1246 50 1318
rect 14 1207 18 1239
rect 70 1208 74 1240
rect 78 1112 82 1320
rect 78 1032 82 1108
rect 126 1112 130 1113
rect -29 164 -25 591
rect -22 274 -18 701
rect -15 384 -11 811
rect -8 494 -4 921
rect -1 604 3 1031
rect 110 1026 114 1100
rect 78 988 82 1018
rect 126 922 130 1108
rect 134 988 138 1018
rect 158 916 162 992
rect 126 878 130 909
rect 182 878 186 913
rect -1 54 3 481
<< m3contact >>
rect -2 1524 2 1528
rect 14 1524 18 1528
rect -28 1515 -24 1519
rect -1 1515 3 1519
rect -29 1141 -25 1145
rect -47 1030 -43 1034
rect -47 920 -43 924
rect -47 810 -43 814
rect 14 1320 18 1324
rect 78 1320 82 1324
rect 14 1239 18 1243
rect 30 1239 34 1243
rect 30 1204 34 1208
rect 70 1204 74 1208
rect 78 1108 82 1112
rect -1 1031 3 1035
rect 126 1108 130 1112
rect -8 921 -4 925
rect -15 811 -11 815
rect -22 701 -18 705
rect -29 591 -25 595
rect 78 1018 82 1022
rect 94 1018 98 1022
rect 94 984 98 988
rect 134 984 138 988
rect 126 909 130 913
rect 142 909 146 913
rect 142 874 146 878
rect 182 874 186 878
rect -1 481 3 485
<< metal3 >>
rect -3 1528 19 1529
rect -3 1524 -2 1528
rect 2 1524 14 1528
rect 18 1524 19 1528
rect -3 1523 19 1524
rect -29 1519 4 1520
rect -29 1515 -28 1519
rect -24 1515 -1 1519
rect 3 1515 4 1519
rect -29 1514 4 1515
rect 13 1324 83 1325
rect 13 1320 14 1324
rect 18 1320 78 1324
rect 82 1320 83 1324
rect 13 1319 83 1320
rect 13 1243 35 1244
rect 13 1239 14 1243
rect 18 1239 30 1243
rect 34 1239 35 1243
rect 13 1238 35 1239
rect 29 1208 75 1209
rect 29 1204 30 1208
rect 34 1204 70 1208
rect 74 1204 75 1208
rect 29 1203 75 1204
rect -30 1145 1 1146
rect -30 1141 -29 1145
rect -25 1141 1 1145
rect -30 1140 1 1141
rect 77 1112 131 1113
rect 77 1108 78 1112
rect 82 1108 126 1112
rect 130 1108 131 1112
rect 77 1107 131 1108
rect -48 1035 0 1036
rect -48 1034 -1 1035
rect -48 1030 -47 1034
rect -43 1031 -1 1034
rect -43 1030 0 1031
rect -48 1029 0 1030
rect 77 1022 99 1023
rect 77 1018 78 1022
rect 82 1018 94 1022
rect 98 1018 99 1022
rect 77 1017 99 1018
rect 93 988 139 989
rect 93 984 94 988
rect 98 984 134 988
rect 138 984 139 988
rect 93 983 139 984
rect -48 925 0 926
rect -48 924 -8 925
rect -48 920 -47 924
rect -43 921 -8 924
rect -4 921 0 925
rect -43 920 0 921
rect -48 919 0 920
rect 125 913 147 914
rect 125 909 126 913
rect 130 909 142 913
rect 146 909 147 913
rect 125 908 147 909
rect 141 878 187 879
rect 141 874 142 878
rect 146 874 182 878
rect 186 874 187 878
rect 141 873 187 874
rect -48 815 0 816
rect -48 814 -15 815
rect -48 810 -47 814
rect -43 811 -15 814
rect -11 811 0 815
rect -43 810 0 811
rect -48 809 0 810
rect -28 705 1 706
rect -28 701 -22 705
rect -18 701 1 705
rect -28 700 1 701
rect -27 595 2 596
rect -25 591 2 595
rect -27 590 2 591
rect -28 485 1 486
rect -28 481 -1 485
rect -28 480 1 481
rect -28 370 1 376
rect -29 260 0 266
rect -28 150 1 156
rect -28 40 1 46
use xor2_2x  xor2_2x_0
timestamp 1492457336
transform 1 0 6 0 1 1214
box -6 -4 74 96
use xor2_2x  xor2_2x_1
timestamp 1492457336
transform 1 0 70 0 1 994
box -6 -4 74 96
use shift_source_gen  shift_source_gen_0
timestamp 1492473219
transform 1 0 -74 0 1 0
box -98 0 162 1648
use xor2_2x  xor2_2x_2
timestamp 1492457336
transform 1 0 118 0 1 884
box -6 -4 74 96
use log_shifter  log_shifter_0
timestamp 1492474365
transform 1 0 112 0 1 0
box -112 0 57 1208
<< labels >>
rlabel metal2 48 1316 48 1316 1 s2
rlabel metal2 112 1098 112 1098 1 s1
rlabel space 64 924 71 926 1 s0
rlabel metal2 160 990 160 990 1 s0
<< end >>
