magic
tech scmos
timestamp 1493746172
<< metal1 >>
rect 30 925 554 940
rect 55 900 529 915
rect 55 887 529 893
rect 195 867 205 870
rect 114 857 119 861
rect 186 848 190 857
rect 131 838 141 841
rect 218 798 253 801
rect 30 787 554 793
rect 445 778 454 782
rect 130 718 134 727
rect 218 723 222 732
rect 226 728 230 737
rect 314 731 317 736
rect 298 728 317 731
rect 266 718 270 727
rect 298 723 302 728
rect 338 723 342 732
rect 377 723 382 732
rect 442 728 446 737
rect 314 720 325 723
rect 250 709 261 712
rect 331 698 342 702
rect 55 687 529 693
rect 419 661 429 664
rect 91 651 101 654
rect 106 648 119 653
rect 322 648 326 657
rect 410 651 414 657
rect 410 648 421 651
rect 298 641 302 647
rect 387 645 397 648
rect 306 641 317 642
rect 298 639 317 641
rect 298 638 309 639
rect 98 631 113 634
rect 298 632 302 638
rect 30 587 554 593
rect 293 578 302 582
rect 375 544 382 552
rect 370 533 413 536
rect 138 518 142 527
rect 290 518 293 533
rect 426 518 430 527
rect 307 515 341 518
rect 250 498 277 501
rect 55 487 529 493
rect 252 478 262 482
rect 178 448 182 459
rect 330 453 334 462
rect 193 448 206 453
rect 158 441 173 444
rect 226 438 237 441
rect 127 428 134 436
rect 226 431 229 438
rect 218 428 229 431
rect 402 398 413 401
rect 30 387 554 393
rect 178 338 182 348
rect 223 344 230 352
rect 186 328 190 337
rect 186 325 205 328
rect 217 323 222 332
rect 346 331 350 337
rect 258 326 269 329
rect 346 328 365 331
rect 418 328 422 337
rect 402 321 406 322
rect 234 318 253 321
rect 387 318 406 321
rect 402 313 406 318
rect 322 310 333 313
rect 55 287 529 293
rect 242 278 253 281
rect 293 278 302 282
rect 410 261 414 264
rect 410 258 421 261
rect 203 247 213 250
rect 266 248 270 257
rect 307 251 325 254
rect 378 248 382 257
rect 138 242 157 245
rect 98 232 102 242
rect 210 238 221 241
rect 418 228 429 231
rect 397 198 406 202
rect 30 187 554 193
rect 258 178 267 182
rect 162 143 166 152
rect 335 144 342 152
rect 378 148 389 151
rect 178 133 182 142
rect 186 138 197 141
rect 194 131 197 138
rect 194 128 205 131
rect 266 128 270 137
rect 115 125 125 128
rect 354 125 365 128
rect 55 87 529 93
rect 55 65 529 80
rect 30 40 554 55
rect 266 28 501 31
<< metal2 >>
rect 18 977 45 980
rect 10 868 13 931
rect 18 848 21 977
rect 30 40 45 940
rect 66 928 69 980
rect 55 65 70 915
rect 98 651 101 980
rect 130 977 141 980
rect 114 858 117 881
rect 106 455 109 651
rect 114 641 117 731
rect 130 721 133 921
rect 138 868 141 977
rect 170 878 173 980
rect 202 867 205 980
rect 322 977 333 980
rect 322 881 325 977
rect 314 878 325 881
rect 146 848 157 851
rect 138 734 141 801
rect 130 718 141 721
rect 114 638 125 641
rect 130 611 133 654
rect 122 608 133 611
rect 82 321 85 454
rect 114 447 117 471
rect 122 428 125 608
rect 138 518 141 718
rect 146 651 149 848
rect 258 828 261 854
rect 274 851 277 861
rect 306 808 309 854
rect 162 748 165 801
rect 234 798 269 801
rect 218 728 221 751
rect 234 721 237 798
rect 290 738 293 801
rect 314 751 317 851
rect 322 838 325 861
rect 330 801 333 844
rect 338 818 341 831
rect 330 798 341 801
rect 314 748 325 751
rect 226 718 237 721
rect 194 698 221 701
rect 162 628 165 641
rect 186 628 189 641
rect 194 621 197 645
rect 202 628 205 661
rect 194 618 205 621
rect 146 478 149 534
rect 130 468 149 471
rect 154 468 157 601
rect 194 598 197 611
rect 186 501 189 521
rect 178 498 189 501
rect 98 331 101 341
rect 82 318 101 321
rect 90 268 93 301
rect 82 198 85 241
rect 98 238 101 318
rect 106 258 109 311
rect 106 58 109 101
rect 114 78 117 421
rect 130 358 133 431
rect 138 418 141 464
rect 146 459 149 468
rect 146 456 157 459
rect 122 331 125 341
rect 138 268 141 312
rect 146 308 149 321
rect 154 319 157 351
rect 162 301 165 461
rect 170 408 173 444
rect 178 418 181 498
rect 146 298 165 301
rect 170 322 173 341
rect 178 338 181 361
rect 186 328 189 341
rect 170 313 174 322
rect 122 248 125 262
rect 122 125 125 151
rect 130 127 133 201
rect 146 168 149 298
rect 154 238 157 271
rect 162 238 165 254
rect 170 228 173 313
rect 194 218 197 521
rect 202 488 205 618
rect 218 551 221 698
rect 226 628 229 718
rect 242 691 245 737
rect 234 688 245 691
rect 234 658 237 688
rect 250 661 253 712
rect 258 678 261 701
rect 282 655 285 671
rect 234 608 237 654
rect 226 598 237 601
rect 218 548 229 551
rect 234 548 237 598
rect 170 128 173 151
rect 178 138 181 161
rect 194 128 197 171
rect 130 118 134 127
rect 170 0 173 111
rect 202 0 205 361
rect 218 348 221 541
rect 226 511 229 548
rect 226 508 237 511
rect 234 471 237 508
rect 226 468 237 471
rect 226 461 229 468
rect 226 381 229 431
rect 242 388 245 445
rect 250 428 253 501
rect 226 378 253 381
rect 210 321 213 332
rect 210 318 221 321
rect 226 318 229 351
rect 234 318 237 351
rect 210 247 213 301
rect 218 281 221 318
rect 242 288 245 334
rect 218 278 245 281
rect 234 231 237 256
rect 210 136 213 231
rect 234 228 245 231
rect 250 228 253 378
rect 258 326 261 361
rect 266 321 269 642
rect 274 578 277 644
rect 290 608 293 734
rect 306 717 309 741
rect 314 708 317 723
rect 322 638 325 748
rect 330 668 333 751
rect 338 728 341 798
rect 346 748 349 801
rect 386 781 389 831
rect 386 778 415 781
rect 346 708 349 734
rect 370 729 373 741
rect 338 661 341 701
rect 330 658 341 661
rect 330 631 333 658
rect 298 578 301 631
rect 314 628 333 631
rect 282 521 285 528
rect 282 518 293 521
rect 306 478 309 521
rect 314 438 317 628
rect 322 548 325 611
rect 338 561 341 653
rect 346 628 349 644
rect 338 558 349 561
rect 330 458 333 531
rect 338 515 341 541
rect 306 351 309 391
rect 338 361 341 401
rect 346 371 349 558
rect 362 541 365 681
rect 370 678 373 711
rect 386 551 389 744
rect 394 645 397 721
rect 402 698 405 771
rect 426 741 429 811
rect 450 778 453 821
rect 410 738 429 741
rect 402 645 405 691
rect 386 548 397 551
rect 362 538 381 541
rect 354 508 357 524
rect 362 518 365 532
rect 346 368 357 371
rect 330 358 341 361
rect 306 348 317 351
rect 266 318 277 321
rect 258 298 261 312
rect 274 298 277 318
rect 282 268 285 324
rect 290 318 293 332
rect 298 278 301 331
rect 306 318 309 332
rect 314 328 317 348
rect 330 331 333 358
rect 330 328 349 331
rect 226 128 230 137
rect 234 125 237 221
rect 242 158 245 228
rect 258 178 261 241
rect 266 188 269 251
rect 290 228 293 241
rect 250 117 253 171
rect 298 115 301 171
rect 234 0 237 111
rect 306 108 309 311
rect 322 268 325 313
rect 322 228 325 254
rect 330 231 333 328
rect 338 298 341 321
rect 338 241 341 271
rect 354 268 357 368
rect 378 341 381 538
rect 394 411 397 548
rect 394 408 405 411
rect 402 361 405 408
rect 362 338 381 341
rect 394 358 405 361
rect 362 315 365 331
rect 370 328 373 338
rect 378 288 381 323
rect 330 228 341 231
rect 338 221 341 228
rect 338 218 349 221
rect 314 125 317 141
rect 346 128 349 218
rect 354 125 357 201
rect 370 198 373 251
rect 378 248 381 271
rect 394 261 397 358
rect 402 318 405 351
rect 410 328 413 738
rect 426 728 445 731
rect 426 678 429 728
rect 434 678 437 701
rect 458 688 461 712
rect 426 541 429 664
rect 426 538 437 541
rect 426 518 429 531
rect 386 258 397 261
rect 386 168 389 258
rect 394 239 397 251
rect 410 231 413 301
rect 418 298 421 491
rect 434 488 437 538
rect 442 518 445 654
rect 410 228 421 231
rect 426 211 429 411
rect 434 288 437 341
rect 442 332 446 342
rect 450 318 453 351
rect 498 301 501 921
rect 490 298 501 301
rect 442 253 445 271
rect 426 208 437 211
rect 402 138 405 201
rect 434 198 437 208
rect 402 135 413 138
rect 450 125 453 191
rect 266 0 269 31
rect 330 0 333 101
rect 338 88 341 101
rect 386 98 389 112
rect 370 0 373 91
rect 402 0 405 124
rect 458 58 461 101
rect 498 28 501 298
rect 514 65 529 915
rect 539 40 554 940
<< metal3 >>
rect 9 927 70 932
rect 0 917 134 922
rect 497 917 584 922
rect 113 877 174 882
rect 9 867 110 872
rect 137 867 278 872
rect 273 862 278 867
rect 273 857 326 862
rect 17 847 150 852
rect 185 847 318 852
rect 137 837 182 842
rect 257 827 390 832
rect 337 817 454 822
rect 305 807 430 812
rect 137 797 222 802
rect 337 767 406 772
rect 161 747 222 752
rect 329 747 350 752
rect 273 737 374 742
rect 113 727 214 732
rect 225 727 366 732
rect 377 727 422 732
rect 265 717 398 722
rect 313 702 318 712
rect 345 707 374 712
rect 257 697 318 702
rect 401 697 438 702
rect 241 687 462 692
rect 361 677 430 682
rect 97 667 254 672
rect 281 667 334 672
rect 249 662 254 667
rect 145 657 238 662
rect 249 657 302 662
rect 377 647 422 652
rect 81 637 126 642
rect 161 637 326 642
rect 97 627 230 632
rect 297 627 350 632
rect 193 607 294 612
rect 241 577 278 582
rect 321 547 382 552
rect 337 537 478 542
rect 137 527 430 532
rect 185 517 286 522
rect 305 517 446 522
rect 353 507 398 512
rect 201 487 254 492
rect 417 487 438 492
rect 257 477 310 482
rect 113 467 158 472
rect 161 457 230 462
rect 201 447 334 452
rect 89 437 190 442
rect 201 437 318 442
rect 121 427 230 432
rect 113 417 182 422
rect 169 407 430 412
rect 337 397 398 402
rect 241 387 310 392
rect 129 357 262 362
rect 153 347 238 352
rect 313 347 406 352
rect 97 337 174 342
rect 185 337 366 342
rect 417 337 446 342
rect 0 327 222 332
rect 257 327 414 332
rect 457 327 486 332
rect 257 322 262 327
rect 145 317 174 322
rect 225 317 262 322
rect 273 317 294 322
rect 305 312 310 322
rect 337 317 454 322
rect 81 307 310 312
rect 0 297 134 302
rect 209 297 422 302
rect 193 287 438 292
rect 0 267 94 272
rect 137 267 158 272
rect 249 267 342 272
rect 353 267 446 272
rect 89 257 374 262
rect 393 257 422 262
rect 369 252 374 257
rect 105 247 230 252
rect 361 247 398 252
rect 81 237 102 242
rect 161 237 294 242
rect 0 227 134 232
rect 169 227 214 232
rect 321 227 414 232
rect 193 217 238 222
rect 0 197 86 202
rect 129 197 190 202
rect 433 192 438 202
rect 241 187 270 192
rect 433 187 454 192
rect 0 167 94 172
rect 145 167 254 172
rect 297 167 390 172
rect 177 157 289 162
rect 121 147 166 152
rect 233 147 286 152
rect 337 147 382 152
rect 281 142 286 147
rect 281 137 318 142
rect 0 127 142 132
rect 169 127 350 132
rect 97 117 134 122
rect 169 107 214 112
rect 233 107 310 112
rect 329 97 390 102
rect 337 87 374 92
rect 0 77 118 82
rect 0 57 110 62
rect 457 57 584 62
use $$M3_M2  $$M3_M2_0
timestamp 1493745683
transform 1 0 12 0 1 930
box -3 -3 3 3
use $$M2_M1_1500_1500_3_3  $$M2_M1_1500_1500_3_3_0
timestamp 1493745683
transform 1 0 37 0 1 932
box -7 -7 7 7
use $$M3_M2  $$M3_M2_1
timestamp 1493745683
transform 1 0 68 0 1 930
box -3 -3 3 3
use $$M2_M1_1500_1500_3_3  $$M2_M1_1500_1500_3_3_1
timestamp 1493745683
transform 1 0 546 0 1 932
box -7 -7 7 7
use $$M3_M2  $$M3_M2_2
timestamp 1493745683
transform 1 0 132 0 1 920
box -3 -3 3 3
use $$M3_M2  $$M3_M2_3
timestamp 1493745683
transform 1 0 500 0 1 920
box -3 -3 3 3
use $$M2_M1_1500_1500_3_3  $$M2_M1_1500_1500_3_3_2
timestamp 1493745683
transform 1 0 62 0 1 907
box -7 -7 7 7
use $$M2_M1_1500_1500_3_3  $$M2_M1_1500_1500_3_3_3
timestamp 1493745683
transform 1 0 521 0 1 907
box -7 -7 7 7
use $$M2_M1_1500_1500_3_1  $$M2_M1_1500_1500_3_1_0
timestamp 1493745683
transform 1 0 62 0 1 890
box -7 -2 7 2
use $$M3_M2  $$M3_M2_5
timestamp 1493745683
transform 1 0 12 0 1 870
box -3 -3 3 3
use $$M3_M2  $$M3_M2_8
timestamp 1493745683
transform 1 0 20 0 1 850
box -3 -3 3 3
use $$M3_M2  $$M3_M2_4
timestamp 1493745683
transform 1 0 116 0 1 880
box -3 -3 3 3
use $$M2_M1  $$M2_M1_0
timestamp 1493745683
transform 1 0 108 0 1 869
box -2 -2 2 2
use $$M3_M2  $$M3_M2_6
timestamp 1493745683
transform 1 0 108 0 1 870
box -3 -3 3 3
use $$M2_M1  $$M2_M1_1
timestamp 1493745683
transform 1 0 116 0 1 860
box -2 -2 2 2
use $$M3_M2  $$M3_M2_7
timestamp 1493745683
transform 1 0 140 0 1 870
box -3 -3 3 3
use $$M2_M1  $$M2_M1_2
timestamp 1493745683
transform 1 0 140 0 1 840
box -2 -2 2 2
use $$M3_M2  $$M3_M2_9
timestamp 1493745683
transform 1 0 140 0 1 840
box -3 -3 3 3
use $$M3_M2  $$M3_M2_10
timestamp 1493745683
transform 1 0 140 0 1 800
box -3 -3 3 3
use $$M3_M2  $$M3_M2_12
timestamp 1493745683
transform 1 0 148 0 1 850
box -3 -3 3 3
use $$M2_M1  $$M2_M1_3
timestamp 1493745683
transform 1 0 156 0 1 853
box -2 -2 2 2
use $$M3_M2  $$M3_M2_11
timestamp 1493745683
transform 1 0 172 0 1 880
box -3 -3 3 3
use $$M2_M1  $$M2_M1_6
timestamp 1493745683
transform 1 0 188 0 1 850
box -2 -2 2 2
use $$M3_M2  $$M3_M2_13
timestamp 1493745683
transform 1 0 188 0 1 850
box -3 -3 3 3
use $$M2_M1  $$M2_M1_7
timestamp 1493745683
transform 1 0 180 0 1 841
box -2 -2 2 2
use $$M3_M2  $$M3_M2_14
timestamp 1493745683
transform 1 0 180 0 1 840
box -3 -3 3 3
use $$M2_M1  $$M2_M1_4
timestamp 1493745683
transform 1 0 164 0 1 800
box -2 -2 2 2
use $$M2_M1  $$M2_M1_5
timestamp 1493745683
transform 1 0 204 0 1 869
box -2 -2 2 2
use $$M2_M1  $$M2_M1_8
timestamp 1493745683
transform 1 0 220 0 1 800
box -2 -2 2 2
use $$M3_M2  $$M3_M2_15
timestamp 1493745683
transform 1 0 220 0 1 800
box -3 -3 3 3
use $$M2_M1  $$M2_M1_9
timestamp 1493745683
transform 1 0 260 0 1 853
box -2 -2 2 2
use $$M3_M2  $$M3_M2_17
timestamp 1493745683
transform 1 0 260 0 1 830
box -3 -3 3 3
use $$M2_M1  $$M2_M1_11
timestamp 1493745683
transform 1 0 268 0 1 800
box -2 -2 2 2
use $$M3_M2  $$M3_M2_16
timestamp 1493745683
transform 1 0 276 0 1 860
box -3 -3 3 3
use $$M2_M1  $$M2_M1_10
timestamp 1493745683
transform 1 0 276 0 1 853
box -2 -2 2 2
use $$M2_M1  $$M2_M1_14
timestamp 1493745683
transform 1 0 292 0 1 800
box -2 -2 2 2
use $$M2_M1  $$M2_M1_12
timestamp 1493745683
transform 1 0 300 0 1 853
box -2 -2 2 2
use $$M2_M1  $$M2_M1_13
timestamp 1493745683
transform 1 0 308 0 1 853
box -2 -2 2 2
use $$M3_M2  $$M3_M2_18
timestamp 1493745683
transform 1 0 300 0 1 850
box -3 -3 3 3
use $$M3_M2  $$M3_M2_19
timestamp 1493745683
transform 1 0 308 0 1 810
box -3 -3 3 3
use $$M2_M1  $$M2_M1_15
timestamp 1493745683
transform 1 0 316 0 1 880
box -2 -2 2 2
use $$M3_M2  $$M3_M2_20
timestamp 1493745683
transform 1 0 324 0 1 860
box -3 -3 3 3
use $$M3_M2  $$M3_M2_21
timestamp 1493745683
transform 1 0 316 0 1 850
box -3 -3 3 3
use $$M2_M1  $$M2_M1_17
timestamp 1493745683
transform 1 0 324 0 1 840
box -2 -2 2 2
use $$M2_M1  $$M2_M1_16
timestamp 1493745683
transform 1 0 332 0 1 843
box -2 -2 2 2
use $$M2_M1  $$M2_M1_18
timestamp 1493745683
transform 1 0 340 0 1 830
box -2 -2 2 2
use $$M3_M2  $$M3_M2_23
timestamp 1493745683
transform 1 0 340 0 1 820
box -3 -3 3 3
use $$M2_M1  $$M2_M1_19
timestamp 1493745683
transform 1 0 348 0 1 800
box -2 -2 2 2
use $$M3_M2  $$M3_M2_22
timestamp 1493745683
transform 1 0 388 0 1 830
box -3 -3 3 3
use $$M3_M2  $$M3_M2_25
timestamp 1493745683
transform 1 0 428 0 1 810
box -3 -3 3 3
use $$M3_M2  $$M3_M2_24
timestamp 1493745683
transform 1 0 452 0 1 820
box -3 -3 3 3
use $$M2_M1_1500_1500_3_1  $$M2_M1_1500_1500_3_1_1
timestamp 1493745683
transform 1 0 521 0 1 890
box -7 -2 7 2
use $$M2_M1_1500_1500_3_1  $$M2_M1_1500_1500_3_1_2
timestamp 1493745683
transform 1 0 37 0 1 790
box -7 -2 7 2
use FILL  FILL_0
timestamp 1493745683
transform 1 0 80 0 -1 890
box -8 -3 16 105
use FILL  FILL_1
timestamp 1493745683
transform 1 0 88 0 -1 890
box -8 -3 16 105
use FILL  FILL_2
timestamp 1493745683
transform 1 0 96 0 -1 890
box -8 -3 16 105
use OR2X1  OR2X1_0
timestamp 1493745683
transform 1 0 104 0 -1 890
box -8 -3 40 105
use FILL  FILL_3
timestamp 1493745683
transform 1 0 136 0 -1 890
box -8 -3 16 105
use FILL  FILL_4
timestamp 1493745683
transform 1 0 144 0 -1 890
box -8 -3 16 105
use INVX2  INVX2_0
timestamp 1493745683
transform 1 0 152 0 -1 890
box -9 -3 26 105
use FILL  FILL_5
timestamp 1493745683
transform 1 0 168 0 -1 890
box -8 -3 16 105
use NOR2X1  NOR2X1_0
timestamp 1493745683
transform -1 0 200 0 -1 890
box -8 -3 32 105
use FILL  FILL_6
timestamp 1493745683
transform 1 0 200 0 -1 890
box -8 -3 16 105
use FILL  FILL_7
timestamp 1493745683
transform 1 0 208 0 -1 890
box -8 -3 16 105
use FILL  FILL_8
timestamp 1493745683
transform 1 0 216 0 -1 890
box -8 -3 16 105
use FILL  FILL_9
timestamp 1493745683
transform 1 0 224 0 -1 890
box -8 -3 16 105
use FILL  FILL_10
timestamp 1493745683
transform 1 0 232 0 -1 890
box -8 -3 16 105
use FILL  FILL_11
timestamp 1493745683
transform 1 0 240 0 -1 890
box -8 -3 16 105
use INVX2  INVX2_1
timestamp 1493745683
transform -1 0 264 0 -1 890
box -9 -3 26 105
use INVX2  INVX2_2
timestamp 1493745683
transform -1 0 280 0 -1 890
box -9 -3 26 105
use FILL  FILL_12
timestamp 1493745683
transform 1 0 280 0 -1 890
box -8 -3 16 105
use INVX2  INVX2_3
timestamp 1493745683
transform -1 0 304 0 -1 890
box -9 -3 26 105
use INVX2  INVX2_4
timestamp 1493745683
transform 1 0 304 0 -1 890
box -9 -3 26 105
use NAND3X1  NAND3X1_0
timestamp 1493745683
transform 1 0 320 0 -1 890
box -8 -3 40 105
use FILL  FILL_13
timestamp 1493745683
transform 1 0 352 0 -1 890
box -8 -3 16 105
use FILL  FILL_14
timestamp 1493745683
transform 1 0 360 0 -1 890
box -8 -3 16 105
use FILL  FILL_15
timestamp 1493745683
transform 1 0 368 0 -1 890
box -8 -3 16 105
use FILL  FILL_16
timestamp 1493745683
transform 1 0 376 0 -1 890
box -8 -3 16 105
use FILL  FILL_17
timestamp 1493745683
transform 1 0 384 0 -1 890
box -8 -3 16 105
use FILL  FILL_18
timestamp 1493745683
transform 1 0 392 0 -1 890
box -8 -3 16 105
use FILL  FILL_19
timestamp 1493745683
transform 1 0 400 0 -1 890
box -8 -3 16 105
use FILL  FILL_20
timestamp 1493745683
transform 1 0 408 0 -1 890
box -8 -3 16 105
use FILL  FILL_21
timestamp 1493745683
transform 1 0 416 0 -1 890
box -8 -3 16 105
use FILL  FILL_22
timestamp 1493745683
transform 1 0 424 0 -1 890
box -8 -3 16 105
use FILL  FILL_23
timestamp 1493745683
transform 1 0 432 0 -1 890
box -8 -3 16 105
use FILL  FILL_24
timestamp 1493745683
transform 1 0 440 0 -1 890
box -8 -3 16 105
use FILL  FILL_25
timestamp 1493745683
transform 1 0 448 0 -1 890
box -8 -3 16 105
use FILL  FILL_26
timestamp 1493745683
transform 1 0 456 0 -1 890
box -8 -3 16 105
use FILL  FILL_27
timestamp 1493745683
transform 1 0 464 0 -1 890
box -8 -3 16 105
use FILL  FILL_28
timestamp 1493745683
transform 1 0 472 0 -1 890
box -8 -3 16 105
use FILL  FILL_29
timestamp 1493745683
transform 1 0 480 0 -1 890
box -8 -3 16 105
use FILL  FILL_30
timestamp 1493745683
transform 1 0 488 0 -1 890
box -8 -3 16 105
use FILL  FILL_31
timestamp 1493745683
transform 1 0 496 0 -1 890
box -8 -3 16 105
use $$M2_M1_1500_1500_3_1  $$M2_M1_1500_1500_3_1_3
timestamp 1493745683
transform 1 0 546 0 1 790
box -7 -2 7 2
use $$M3_M2  $$M3_M2_26
timestamp 1493745683
transform 1 0 164 0 1 750
box -3 -3 3 3
use $$M2_M1  $$M2_M1_20
timestamp 1493745683
transform 1 0 140 0 1 736
box -2 -2 2 2
use $$M3_M2  $$M3_M2_27
timestamp 1493745683
transform 1 0 116 0 1 730
box -3 -3 3 3
use $$M2_M1  $$M2_M1_21
timestamp 1493745683
transform 1 0 132 0 1 720
box -2 -2 2 2
use $$M2_M1  $$M2_M1_22
timestamp 1493745683
transform 1 0 196 0 1 700
box -2 -2 2 2
use $$M3_M2  $$M3_M2_28
timestamp 1493745683
transform 1 0 220 0 1 750
box -3 -3 3 3
use $$M2_M1  $$M2_M1_23
timestamp 1493745683
transform 1 0 244 0 1 736
box -2 -2 2 2
use $$M2_M1  $$M2_M1_24
timestamp 1493745683
transform 1 0 212 0 1 733
box -2 -2 2 2
use $$M3_M2  $$M3_M2_29
timestamp 1493745683
transform 1 0 212 0 1 730
box -3 -3 3 3
use $$M2_M1  $$M2_M1_25
timestamp 1493745683
transform 1 0 220 0 1 730
box -2 -2 2 2
use $$M2_M1  $$M2_M1_26
timestamp 1493745683
transform 1 0 228 0 1 730
box -2 -2 2 2
use $$M3_M2  $$M3_M2_30
timestamp 1493745683
transform 1 0 228 0 1 730
box -3 -3 3 3
use $$M2_M1  $$M2_M1_27
timestamp 1493745683
transform 1 0 236 0 1 724
box -2 -2 2 2
use $$M2_M1  $$M2_M1_30
timestamp 1493745683
transform 1 0 252 0 1 711
box -2 -2 2 2
use $$M2_M1  $$M2_M1_28
timestamp 1493745683
transform 1 0 276 0 1 739
box -2 -2 2 2
use $$M3_M2  $$M3_M2_31
timestamp 1493745683
transform 1 0 276 0 1 740
box -3 -3 3 3
use $$M2_M1  $$M2_M1_29
timestamp 1493745683
transform 1 0 268 0 1 720
box -2 -2 2 2
use $$M3_M2  $$M3_M2_32
timestamp 1493745683
transform 1 0 268 0 1 720
box -3 -3 3 3
use $$M3_M2  $$M3_M2_33
timestamp 1493745683
transform 1 0 260 0 1 700
box -3 -3 3 3
use $$M3_M2  $$M3_M2_37
timestamp 1493745683
transform 1 0 292 0 1 740
box -3 -3 3 3
use $$M2_M1  $$M2_M1_31
timestamp 1493745683
transform 1 0 292 0 1 733
box -2 -2 2 2
use $$M3_M2  $$M3_M2_34
timestamp 1493745683
transform 1 0 340 0 1 770
box -3 -3 3 3
use $$M3_M2  $$M3_M2_35
timestamp 1493745683
transform 1 0 332 0 1 750
box -3 -3 3 3
use $$M3_M2  $$M3_M2_36
timestamp 1493745683
transform 1 0 348 0 1 750
box -3 -3 3 3
use $$M3_M2  $$M3_M2_38
timestamp 1493745683
transform 1 0 308 0 1 740
box -3 -3 3 3
use $$M2_M1  $$M2_M1_33
timestamp 1493745683
transform 1 0 340 0 1 730
box -2 -2 2 2
use $$M2_M1  $$M2_M1_32
timestamp 1493745683
transform 1 0 348 0 1 733
box -2 -2 2 2
use $$M2_M1  $$M2_M1_35
timestamp 1493745683
transform 1 0 308 0 1 718
box -2 -2 2 2
use $$M2_M1  $$M2_M1_34
timestamp 1493745683
transform 1 0 316 0 1 721
box -2 -2 2 2
use $$M3_M2  $$M3_M2_39
timestamp 1493745683
transform 1 0 316 0 1 710
box -3 -3 3 3
use $$M3_M2  $$M3_M2_40
timestamp 1493745683
transform 1 0 348 0 1 710
box -3 -3 3 3
use $$M2_M1  $$M2_M1_36
timestamp 1493745683
transform 1 0 340 0 1 700
box -2 -2 2 2
use $$M3_M2  $$M3_M2_41
timestamp 1493745683
transform 1 0 372 0 1 740
box -3 -3 3 3
use $$M2_M1  $$M2_M1_37
timestamp 1493745683
transform 1 0 388 0 1 743
box -2 -2 2 2
use $$M3_M2  $$M3_M2_42
timestamp 1493745683
transform 1 0 364 0 1 730
box -3 -3 3 3
use $$M2_M1  $$M2_M1_38
timestamp 1493745683
transform 1 0 372 0 1 731
box -2 -2 2 2
use $$M2_M1  $$M2_M1_39
timestamp 1493745683
transform 1 0 380 0 1 730
box -2 -2 2 2
use $$M3_M2  $$M3_M2_43
timestamp 1493745683
transform 1 0 380 0 1 730
box -3 -3 3 3
use $$M2_M1  $$M2_M1_40
timestamp 1493745683
transform 1 0 364 0 1 727
box -2 -2 2 2
use $$M2_M1  $$M2_M1_41
timestamp 1493745683
transform 1 0 414 0 1 780
box -2 -2 2 2
use $$M3_M2  $$M3_M2_44
timestamp 1493745683
transform 1 0 404 0 1 770
box -3 -3 3 3
use $$M2_M1  $$M2_M1_42
timestamp 1493745683
transform 1 0 404 0 1 744
box -2 -2 2 2
use $$M2_M1  $$M2_M1_43
timestamp 1493745683
transform 1 0 420 0 1 731
box -2 -2 2 2
use $$M3_M2  $$M3_M2_45
timestamp 1493745683
transform 1 0 420 0 1 730
box -3 -3 3 3
use $$M3_M2  $$M3_M2_46
timestamp 1493745683
transform 1 0 396 0 1 720
box -3 -3 3 3
use $$M3_M2  $$M3_M2_47
timestamp 1493745683
transform 1 0 372 0 1 710
box -3 -3 3 3
use $$M3_M2  $$M3_M2_48
timestamp 1493745683
transform 1 0 404 0 1 700
box -3 -3 3 3
use $$M2_M1  $$M2_M1_44
timestamp 1493745683
transform 1 0 428 0 1 727
box -2 -2 2 2
use $$M2_M1  $$M2_M1_45
timestamp 1493745683
transform 1 0 452 0 1 780
box -2 -2 2 2
use $$M2_M1  $$M2_M1_46
timestamp 1493745683
transform 1 0 444 0 1 730
box -2 -2 2 2
use $$M3_M2  $$M3_M2_49
timestamp 1493745683
transform 1 0 436 0 1 700
box -3 -3 3 3
use $$M2_M1  $$M2_M1_47
timestamp 1493745683
transform 1 0 460 0 1 711
box -2 -2 2 2
use $$M2_M1_1500_1500_3_1  $$M2_M1_1500_1500_3_1_4
timestamp 1493745683
transform 1 0 62 0 1 690
box -7 -2 7 2
use FILL  FILL_32
timestamp 1493745683
transform -1 0 88 0 1 690
box -8 -3 16 105
use FILL  FILL_33
timestamp 1493745683
transform -1 0 96 0 1 690
box -8 -3 16 105
use FILL  FILL_34
timestamp 1493745683
transform -1 0 104 0 1 690
box -8 -3 16 105
use DFFPOSX1  DFFPOSX1_0
timestamp 1493147875
transform 1 0 104 0 1 690
box -8 -3 104 105
use FILL  FILL_36
timestamp 1493745683
transform -1 0 208 0 1 690
box -8 -3 16 105
use $$M3_M2  $$M3_M2_50
timestamp 1493745683
transform 1 0 244 0 1 690
box -3 -3 3 3
use AOI22X1  AOI22X1_0
timestamp 1493147875
transform -1 0 248 0 1 690
box -8 -3 46 105
use FILL  FILL_42
timestamp 1493745683
transform -1 0 256 0 1 690
box -8 -3 16 105
use NOR2X1  NOR2X1_1
timestamp 1493745683
transform 1 0 256 0 1 690
box -8 -3 32 105
use FILL  FILL_43
timestamp 1493745683
transform -1 0 288 0 1 690
box -8 -3 16 105
use NOR2X1  NOR2X1_2
timestamp 1493745683
transform -1 0 312 0 1 690
box -8 -3 32 105
use AOI22X1  AOI22X1_1
timestamp 1493147875
transform 1 0 312 0 1 690
box -8 -3 46 105
use FILL  FILL_46
timestamp 1493745683
transform -1 0 360 0 1 690
box -8 -3 16 105
use OAI21X1  OAI21X1_0
timestamp 1493745683
transform 1 0 360 0 1 690
box -8 -3 34 105
use $$M3_M2  $$M3_M2_51
timestamp 1493745683
transform 1 0 404 0 1 690
box -3 -3 3 3
use FILL  FILL_48
timestamp 1493745683
transform -1 0 400 0 1 690
box -8 -3 16 105
use OAI21X1  OAI21X1_1
timestamp 1493745683
transform -1 0 432 0 1 690
box -8 -3 34 105
use FILL  FILL_49
timestamp 1493745683
transform -1 0 440 0 1 690
box -8 -3 16 105
use $$M3_M2  $$M3_M2_52
timestamp 1493745683
transform 1 0 460 0 1 690
box -3 -3 3 3
use NOR2X1  NOR2X1_3
timestamp 1493745683
transform -1 0 464 0 1 690
box -8 -3 32 105
use FILL  FILL_50
timestamp 1493745683
transform -1 0 472 0 1 690
box -8 -3 16 105
use FILL  FILL_51
timestamp 1493745683
transform -1 0 480 0 1 690
box -8 -3 16 105
use FILL  FILL_52
timestamp 1493745683
transform -1 0 488 0 1 690
box -8 -3 16 105
use FILL  FILL_53
timestamp 1493745683
transform -1 0 496 0 1 690
box -8 -3 16 105
use FILL  FILL_54
timestamp 1493745683
transform -1 0 504 0 1 690
box -8 -3 16 105
use $$M2_M1_1500_1500_3_1  $$M2_M1_1500_1500_3_1_5
timestamp 1493745683
transform 1 0 521 0 1 690
box -7 -2 7 2
use $$M3_M2  $$M3_M2_53
timestamp 1493745683
transform 1 0 100 0 1 670
box -3 -3 3 3
use $$M2_M1  $$M2_M1_48
timestamp 1493745683
transform 1 0 100 0 1 653
box -2 -2 2 2
use $$M2_M1  $$M2_M1_49
timestamp 1493745683
transform 1 0 84 0 1 640
box -2 -2 2 2
use $$M3_M2  $$M3_M2_54
timestamp 1493745683
transform 1 0 84 0 1 640
box -3 -3 3 3
use $$M2_M1  $$M2_M1_52
timestamp 1493745683
transform 1 0 108 0 1 650
box -2 -2 2 2
use $$M2_M1  $$M2_M1_50
timestamp 1493745683
transform 1 0 100 0 1 633
box -2 -2 2 2
use $$M3_M2  $$M3_M2_55
timestamp 1493745683
transform 1 0 100 0 1 630
box -3 -3 3 3
use $$M2_M1  $$M2_M1_51
timestamp 1493745683
transform 1 0 132 0 1 653
box -2 -2 2 2
use $$M2_M1  $$M2_M1_53
timestamp 1493745683
transform 1 0 124 0 1 642
box -2 -2 2 2
use $$M3_M2  $$M3_M2_56
timestamp 1493745683
transform 1 0 124 0 1 640
box -3 -3 3 3
use $$M3_M2  $$M3_M2_57
timestamp 1493745683
transform 1 0 148 0 1 660
box -3 -3 3 3
use $$M2_M1  $$M2_M1_54
timestamp 1493745683
transform 1 0 148 0 1 653
box -2 -2 2 2
use $$M3_M2  $$M3_M2_59
timestamp 1493745683
transform 1 0 164 0 1 640
box -3 -3 3 3
use $$M2_M1  $$M2_M1_57
timestamp 1493745683
transform 1 0 164 0 1 630
box -2 -2 2 2
use $$M2_M1  $$M2_M1_59
timestamp 1493745683
transform 1 0 156 0 1 600
box -2 -2 2 2
use $$M3_M2  $$M3_M2_58
timestamp 1493745683
transform 1 0 204 0 1 660
box -3 -3 3 3
use $$M2_M1  $$M2_M1_55
timestamp 1493745683
transform 1 0 196 0 1 644
box -2 -2 2 2
use $$M2_M1  $$M2_M1_56
timestamp 1493745683
transform 1 0 188 0 1 640
box -2 -2 2 2
use $$M3_M2  $$M3_M2_60
timestamp 1493745683
transform 1 0 188 0 1 630
box -3 -3 3 3
use $$M2_M1  $$M2_M1_58
timestamp 1493745683
transform 1 0 204 0 1 630
box -2 -2 2 2
use $$M3_M2  $$M3_M2_61
timestamp 1493745683
transform 1 0 196 0 1 610
box -3 -3 3 3
use $$M2_M1  $$M2_M1_60
timestamp 1493745683
transform 1 0 196 0 1 600
box -2 -2 2 2
use $$M3_M2  $$M3_M2_62
timestamp 1493745683
transform 1 0 236 0 1 660
box -3 -3 3 3
use $$M2_M1  $$M2_M1_61
timestamp 1493745683
transform 1 0 236 0 1 653
box -2 -2 2 2
use $$M3_M2  $$M3_M2_63
timestamp 1493745683
transform 1 0 228 0 1 630
box -3 -3 3 3
use $$M3_M2  $$M3_M2_64
timestamp 1493745683
transform 1 0 236 0 1 610
box -3 -3 3 3
use $$M2_M1  $$M2_M1_62
timestamp 1493745683
transform 1 0 228 0 1 600
box -2 -2 2 2
use $$M2_M1  $$M2_M1_63
timestamp 1493745683
transform 1 0 260 0 1 680
box -2 -2 2 2
use $$M3_M2  $$M3_M2_65
timestamp 1493745683
transform 1 0 252 0 1 670
box -3 -3 3 3
use $$M2_M1  $$M2_M1_64
timestamp 1493745683
transform 1 0 252 0 1 663
box -2 -2 2 2
use $$M3_M2  $$M3_M2_66
timestamp 1493745683
transform 1 0 284 0 1 670
box -3 -3 3 3
use $$M2_M1  $$M2_M1_66
timestamp 1493745683
transform 1 0 284 0 1 657
box -2 -2 2 2
use $$M2_M1  $$M2_M1_65
timestamp 1493745683
transform 1 0 300 0 1 663
box -2 -2 2 2
use $$M3_M2  $$M3_M2_67
timestamp 1493745683
transform 1 0 300 0 1 660
box -3 -3 3 3
use $$M2_M1  $$M2_M1_68
timestamp 1493745683
transform 1 0 268 0 1 641
box -2 -2 2 2
use $$M2_M1  $$M2_M1_67
timestamp 1493745683
transform 1 0 276 0 1 643
box -2 -2 2 2
use $$M3_M2  $$M3_M2_68
timestamp 1493745683
transform 1 0 300 0 1 630
box -3 -3 3 3
use $$M3_M2  $$M3_M2_69
timestamp 1493745683
transform 1 0 292 0 1 610
box -3 -3 3 3
use $$M3_M2  $$M3_M2_70
timestamp 1493745683
transform 1 0 332 0 1 670
box -3 -3 3 3
use $$M2_M1  $$M2_M1_70
timestamp 1493745683
transform 1 0 324 0 1 650
box -2 -2 2 2
use $$M2_M1  $$M2_M1_69
timestamp 1493745683
transform 1 0 340 0 1 652
box -2 -2 2 2
use $$M3_M2  $$M3_M2_71
timestamp 1493745683
transform 1 0 324 0 1 640
box -3 -3 3 3
use $$M2_M1  $$M2_M1_71
timestamp 1493745683
transform 1 0 348 0 1 643
box -2 -2 2 2
use $$M3_M2  $$M3_M2_72
timestamp 1493745683
transform 1 0 348 0 1 630
box -3 -3 3 3
use $$M2_M1  $$M2_M1_72
timestamp 1493745683
transform 1 0 324 0 1 610
box -2 -2 2 2
use $$M3_M2  $$M3_M2_73
timestamp 1493745683
transform 1 0 364 0 1 680
box -3 -3 3 3
use $$M2_M1  $$M2_M1_73
timestamp 1493745683
transform 1 0 372 0 1 680
box -2 -2 2 2
use $$M2_M1  $$M2_M1_74
timestamp 1493745683
transform 1 0 364 0 1 667
box -2 -2 2 2
use $$M2_M1  $$M2_M1_75
timestamp 1493745683
transform 1 0 380 0 1 652
box -2 -2 2 2
use $$M3_M2  $$M3_M2_74
timestamp 1493745683
transform 1 0 380 0 1 650
box -3 -3 3 3
use $$M2_M1  $$M2_M1_79
timestamp 1493745683
transform 1 0 396 0 1 647
box -2 -2 2 2
use $$M2_M1  $$M2_M1_80
timestamp 1493745683
transform 1 0 404 0 1 647
box -2 -2 2 2
use $$M3_M2  $$M3_M2_75
timestamp 1493745683
transform 1 0 428 0 1 680
box -3 -3 3 3
use $$M2_M1  $$M2_M1_76
timestamp 1493745683
transform 1 0 436 0 1 680
box -2 -2 2 2
use $$M2_M1  $$M2_M1_77
timestamp 1493745683
transform 1 0 428 0 1 663
box -2 -2 2 2
use $$M2_M1  $$M2_M1_78
timestamp 1493745683
transform 1 0 420 0 1 650
box -2 -2 2 2
use $$M3_M2  $$M3_M2_76
timestamp 1493745683
transform 1 0 420 0 1 650
box -3 -3 3 3
use $$M2_M1  $$M2_M1_81
timestamp 1493745683
transform 1 0 444 0 1 653
box -2 -2 2 2
use $$M2_M1_1500_1500_3_1  $$M2_M1_1500_1500_3_1_6
timestamp 1493745683
transform 1 0 37 0 1 590
box -7 -2 7 2
use INVX2  INVX2_5
timestamp 1493745683
transform -1 0 96 0 -1 690
box -9 -3 26 105
use FILL  FILL_35
timestamp 1493745683
transform 1 0 96 0 -1 690
box -8 -3 16 105
use OAI21X1  OAI21X1_2
timestamp 1493745683
transform -1 0 136 0 -1 690
box -8 -3 34 105
use FILL  FILL_37
timestamp 1493745683
transform 1 0 136 0 -1 690
box -8 -3 16 105
use NAND2X1  NAND2X1_0
timestamp 1493745683
transform 1 0 144 0 -1 690
box -8 -3 32 105
use FILL  FILL_38
timestamp 1493745683
transform 1 0 168 0 -1 690
box -8 -3 16 105
use FILL  FILL_39
timestamp 1493745683
transform 1 0 176 0 -1 690
box -8 -3 16 105
use NAND3X1  NAND3X1_1
timestamp 1493745683
transform 1 0 184 0 -1 690
box -8 -3 40 105
use FILL  FILL_40
timestamp 1493745683
transform 1 0 216 0 -1 690
box -8 -3 16 105
use INVX2  INVX2_6
timestamp 1493745683
transform -1 0 240 0 -1 690
box -9 -3 26 105
use FILL  FILL_41
timestamp 1493745683
transform 1 0 240 0 -1 690
box -8 -3 16 105
use NOR2X1  NOR2X1_4
timestamp 1493745683
transform 1 0 248 0 -1 690
box -8 -3 32 105
use AOI21X1  AOI21X1_0
timestamp 1493745683
transform 1 0 272 0 -1 690
box -7 -3 39 105
use FILL  FILL_44
timestamp 1493745683
transform 1 0 304 0 -1 690
box -8 -3 16 105
use AOI22X1  AOI22X1_2
timestamp 1493147875
transform -1 0 352 0 -1 690
box -8 -3 46 105
use FILL  FILL_45
timestamp 1493745683
transform 1 0 352 0 -1 690
box -8 -3 16 105
use AOI21X1  AOI21X1_1
timestamp 1493745683
transform -1 0 392 0 -1 690
box -7 -3 39 105
use FILL  FILL_47
timestamp 1493745683
transform 1 0 392 0 -1 690
box -8 -3 16 105
use NOR2X1  NOR2X1_5
timestamp 1493745683
transform -1 0 424 0 -1 690
box -8 -3 32 105
use FILL  FILL_55
timestamp 1493745683
transform 1 0 424 0 -1 690
box -8 -3 16 105
use INVX2  INVX2_7
timestamp 1493745683
transform -1 0 448 0 -1 690
box -9 -3 26 105
use FILL  FILL_56
timestamp 1493745683
transform 1 0 448 0 -1 690
box -8 -3 16 105
use FILL  FILL_57
timestamp 1493745683
transform 1 0 456 0 -1 690
box -8 -3 16 105
use FILL  FILL_58
timestamp 1493745683
transform 1 0 464 0 -1 690
box -8 -3 16 105
use FILL  FILL_59
timestamp 1493745683
transform 1 0 472 0 -1 690
box -8 -3 16 105
use FILL  FILL_60
timestamp 1493745683
transform 1 0 480 0 -1 690
box -8 -3 16 105
use FILL  FILL_61
timestamp 1493745683
transform 1 0 488 0 -1 690
box -8 -3 16 105
use FILL  FILL_62
timestamp 1493745683
transform 1 0 496 0 -1 690
box -8 -3 16 105
use $$M2_M1_1500_1500_3_1  $$M2_M1_1500_1500_3_1_7
timestamp 1493745683
transform 1 0 546 0 1 590
box -7 -2 7 2
use $$M3_M2  $$M3_M2_77
timestamp 1493745683
transform 1 0 140 0 1 530
box -3 -3 3 3
use $$M2_M1  $$M2_M1_82
timestamp 1493745683
transform 1 0 148 0 1 533
box -2 -2 2 2
use $$M2_M1  $$M2_M1_83
timestamp 1493745683
transform 1 0 140 0 1 520
box -2 -2 2 2
use $$M3_M2  $$M3_M2_78
timestamp 1493745683
transform 1 0 188 0 1 520
box -3 -3 3 3
use $$M2_M1  $$M2_M1_84
timestamp 1493745683
transform 1 0 196 0 1 520
box -2 -2 2 2
use $$M2_M1  $$M2_M1_85
timestamp 1493745683
transform 1 0 244 0 1 580
box -2 -2 2 2
use $$M3_M2  $$M3_M2_79
timestamp 1493745683
transform 1 0 244 0 1 580
box -3 -3 3 3
use $$M2_M1  $$M2_M1_86
timestamp 1493745683
transform 1 0 236 0 1 550
box -2 -2 2 2
use $$M2_M1  $$M2_M1_87
timestamp 1493745683
transform 1 0 220 0 1 540
box -2 -2 2 2
use $$M2_M1  $$M2_M1_88
timestamp 1493745683
transform 1 0 228 0 1 534
box -2 -2 2 2
use $$M2_M1  $$M2_M1_89
timestamp 1493745683
transform 1 0 252 0 1 500
box -2 -2 2 2
use $$M3_M2  $$M3_M2_80
timestamp 1493745683
transform 1 0 276 0 1 580
box -3 -3 3 3
use $$M2_M1  $$M2_M1_90
timestamp 1493745683
transform 1 0 300 0 1 580
box -2 -2 2 2
use $$M2_M1  $$M2_M1_91
timestamp 1493745683
transform 1 0 284 0 1 527
box -2 -2 2 2
use $$M3_M2  $$M3_M2_85
timestamp 1493745683
transform 1 0 284 0 1 520
box -3 -3 3 3
use $$M2_M1  $$M2_M1_94
timestamp 1493745683
transform 1 0 292 0 1 520
box -2 -2 2 2
use $$M3_M2  $$M3_M2_86
timestamp 1493745683
transform 1 0 308 0 1 520
box -3 -3 3 3
use $$M3_M2  $$M3_M2_81
timestamp 1493745683
transform 1 0 324 0 1 550
box -3 -3 3 3
use $$M3_M2  $$M3_M2_83
timestamp 1493745683
transform 1 0 340 0 1 540
box -3 -3 3 3
use $$M3_M2  $$M3_M2_84
timestamp 1493745683
transform 1 0 332 0 1 530
box -3 -3 3 3
use $$M2_M1  $$M2_M1_96
timestamp 1493745683
transform 1 0 340 0 1 517
box -2 -2 2 2
use $$M2_M1  $$M2_M1_92
timestamp 1493745683
transform 1 0 380 0 1 550
box -2 -2 2 2
use $$M3_M2  $$M3_M2_82
timestamp 1493745683
transform 1 0 380 0 1 550
box -3 -3 3 3
use $$M2_M1  $$M2_M1_93
timestamp 1493745683
transform 1 0 364 0 1 531
box -2 -2 2 2
use $$M2_M1  $$M2_M1_95
timestamp 1493745683
transform 1 0 356 0 1 523
box -2 -2 2 2
use $$M3_M2  $$M3_M2_87
timestamp 1493745683
transform 1 0 364 0 1 520
box -3 -3 3 3
use $$M3_M2  $$M3_M2_88
timestamp 1493745683
transform 1 0 356 0 1 510
box -3 -3 3 3
use $$M3_M2  $$M3_M2_93
timestamp 1493745683
transform 1 0 396 0 1 510
box -3 -3 3 3
use $$M3_M2  $$M3_M2_89
timestamp 1493745683
transform 1 0 436 0 1 540
box -3 -3 3 3
use $$M2_M1  $$M2_M1_97
timestamp 1493745683
transform 1 0 476 0 1 540
box -2 -2 2 2
use $$M3_M2  $$M3_M2_90
timestamp 1493745683
transform 1 0 476 0 1 540
box -3 -3 3 3
use $$M3_M2  $$M3_M2_91
timestamp 1493745683
transform 1 0 428 0 1 530
box -3 -3 3 3
use $$M2_M1  $$M2_M1_98
timestamp 1493745683
transform 1 0 428 0 1 520
box -2 -2 2 2
use $$M3_M2  $$M3_M2_92
timestamp 1493745683
transform 1 0 444 0 1 520
box -3 -3 3 3
use $$M2_M1_1500_1500_3_1  $$M2_M1_1500_1500_3_1_8
timestamp 1493745683
transform 1 0 62 0 1 490
box -7 -2 7 2
use FILL  FILL_63
timestamp 1493745683
transform -1 0 88 0 1 490
box -8 -3 16 105
use FILL  FILL_64
timestamp 1493745683
transform -1 0 96 0 1 490
box -8 -3 16 105
use FILL  FILL_65
timestamp 1493745683
transform -1 0 104 0 1 490
box -8 -3 16 105
use FILL  FILL_67
timestamp 1493745683
transform -1 0 112 0 1 490
box -8 -3 16 105
use $$M3_M2  $$M3_M2_94
timestamp 1493745683
transform 1 0 204 0 1 490
box -3 -3 3 3
use DFFPOSX1  DFFPOSX1_1
timestamp 1493147875
transform 1 0 112 0 1 490
box -8 -3 104 105
use FILL  FILL_69
timestamp 1493745683
transform -1 0 216 0 1 490
box -8 -3 16 105
use $$M3_M2  $$M3_M2_95
timestamp 1493745683
transform 1 0 252 0 1 490
box -3 -3 3 3
use NAND3X1  NAND3X1_2
timestamp 1493745683
transform 1 0 216 0 1 490
box -8 -3 40 105
use FILL  FILL_71
timestamp 1493745683
transform -1 0 256 0 1 490
box -8 -3 16 105
use FILL  FILL_72
timestamp 1493745683
transform -1 0 264 0 1 490
box -8 -3 16 105
use FILL  FILL_73
timestamp 1493745683
transform -1 0 272 0 1 490
box -8 -3 16 105
use INVX2  INVX2_8
timestamp 1493745683
transform -1 0 288 0 1 490
box -9 -3 26 105
use NOR2X1  NOR2X1_6
timestamp 1493745683
transform -1 0 312 0 1 490
box -8 -3 32 105
use FILL  FILL_74
timestamp 1493745683
transform -1 0 320 0 1 490
box -8 -3 16 105
use FILL  FILL_75
timestamp 1493745683
transform -1 0 328 0 1 490
box -8 -3 16 105
use FILL  FILL_76
timestamp 1493745683
transform -1 0 336 0 1 490
box -8 -3 16 105
use FILL  FILL_77
timestamp 1493745683
transform -1 0 344 0 1 490
box -8 -3 16 105
use FILL  FILL_78
timestamp 1493745683
transform -1 0 352 0 1 490
box -8 -3 16 105
use OAI21X1  OAI21X1_3
timestamp 1493745683
transform 1 0 352 0 1 490
box -8 -3 34 105
use FILL  FILL_79
timestamp 1493745683
transform -1 0 392 0 1 490
box -8 -3 16 105
use FILL  FILL_85
timestamp 1493745683
transform -1 0 400 0 1 490
box -8 -3 16 105
use $$M3_M2  $$M3_M2_96
timestamp 1493745683
transform 1 0 420 0 1 490
box -3 -3 3 3
use $$M3_M2  $$M3_M2_97
timestamp 1493745683
transform 1 0 436 0 1 490
box -3 -3 3 3
use DFFPOSX1  DFFPOSX1_2
timestamp 1493147875
transform 1 0 400 0 1 490
box -8 -3 104 105
use FILL  FILL_86
timestamp 1493745683
transform -1 0 504 0 1 490
box -8 -3 16 105
use $$M2_M1_1500_1500_3_1  $$M2_M1_1500_1500_3_1_9
timestamp 1493745683
transform 1 0 521 0 1 490
box -7 -2 7 2
use $$M2_M1  $$M2_M1_99
timestamp 1493745683
transform 1 0 84 0 1 453
box -2 -2 2 2
use $$M2_M1  $$M2_M1_100
timestamp 1493745683
transform 1 0 92 0 1 440
box -2 -2 2 2
use $$M3_M2  $$M3_M2_98
timestamp 1493745683
transform 1 0 92 0 1 440
box -3 -3 3 3
use $$M3_M2  $$M3_M2_99
timestamp 1493745683
transform 1 0 116 0 1 470
box -3 -3 3 3
use $$M2_M1  $$M2_M1_101
timestamp 1493745683
transform 1 0 148 0 1 480
box -2 -2 2 2
use $$M2_M1  $$M2_M1_102
timestamp 1493745683
transform 1 0 132 0 1 470
box -2 -2 2 2
use $$M2_M1  $$M2_M1_103
timestamp 1493745683
transform 1 0 108 0 1 457
box -2 -2 2 2
use $$M2_M1  $$M2_M1_104
timestamp 1493745683
transform 1 0 116 0 1 449
box -2 -2 2 2
use $$M3_M2  $$M3_M2_102
timestamp 1493745683
transform 1 0 124 0 1 430
box -3 -3 3 3
use $$M3_M2  $$M3_M2_100
timestamp 1493745683
transform 1 0 156 0 1 470
box -3 -3 3 3
use $$M2_M1  $$M2_M1_105
timestamp 1493745683
transform 1 0 140 0 1 463
box -2 -2 2 2
use $$M2_M1  $$M2_M1_106
timestamp 1493745683
transform 1 0 156 0 1 458
box -2 -2 2 2
use $$M3_M2  $$M3_M2_101
timestamp 1493745683
transform 1 0 164 0 1 460
box -3 -3 3 3
use $$M2_M1  $$M2_M1_107
timestamp 1493745683
transform 1 0 132 0 1 430
box -2 -2 2 2
use $$M3_M2  $$M3_M2_103
timestamp 1493745683
transform 1 0 116 0 1 420
box -3 -3 3 3
use $$M3_M2  $$M3_M2_105
timestamp 1493745683
transform 1 0 140 0 1 420
box -3 -3 3 3
use $$M2_M1  $$M2_M1_108
timestamp 1493745683
transform 1 0 180 0 1 450
box -2 -2 2 2
use $$M2_M1  $$M2_M1_110
timestamp 1493745683
transform 1 0 172 0 1 443
box -2 -2 2 2
use $$M2_M1  $$M2_M1_109
timestamp 1493745683
transform 1 0 204 0 1 450
box -2 -2 2 2
use $$M3_M2  $$M3_M2_104
timestamp 1493745683
transform 1 0 204 0 1 450
box -3 -3 3 3
use $$M2_M1  $$M2_M1_111
timestamp 1493745683
transform 1 0 188 0 1 443
box -2 -2 2 2
use $$M3_M2  $$M3_M2_106
timestamp 1493745683
transform 1 0 188 0 1 440
box -3 -3 3 3
use $$M3_M2  $$M3_M2_107
timestamp 1493745683
transform 1 0 204 0 1 440
box -3 -3 3 3
use $$M3_M2  $$M3_M2_108
timestamp 1493745683
transform 1 0 180 0 1 420
box -3 -3 3 3
use $$M3_M2  $$M3_M2_109
timestamp 1493745683
transform 1 0 172 0 1 410
box -3 -3 3 3
use $$M2_M1  $$M2_M1_112
timestamp 1493745683
transform 1 0 204 0 1 437
box -2 -2 2 2
use $$M2_M1  $$M2_M1_114
timestamp 1493745683
transform 1 0 228 0 1 463
box -2 -2 2 2
use $$M3_M2  $$M3_M2_111
timestamp 1493745683
transform 1 0 228 0 1 460
box -3 -3 3 3
use $$M2_M1  $$M2_M1_113
timestamp 1493745683
transform 1 0 260 0 1 480
box -2 -2 2 2
use $$M3_M2  $$M3_M2_110
timestamp 1493745683
transform 1 0 260 0 1 480
box -3 -3 3 3
use $$M2_M1  $$M2_M1_115
timestamp 1493745683
transform 1 0 244 0 1 444
box -2 -2 2 2
use $$M2_M1  $$M2_M1_116
timestamp 1493745683
transform 1 0 228 0 1 430
box -2 -2 2 2
use $$M3_M2  $$M3_M2_112
timestamp 1493745683
transform 1 0 228 0 1 430
box -3 -3 3 3
use $$M2_M1  $$M2_M1_117
timestamp 1493745683
transform 1 0 252 0 1 430
box -2 -2 2 2
use $$M3_M2  $$M3_M2_113
timestamp 1493745683
transform 1 0 308 0 1 480
box -3 -3 3 3
use $$M2_M1  $$M2_M1_118
timestamp 1493745683
transform 1 0 332 0 1 460
box -2 -2 2 2
use $$M3_M2  $$M3_M2_114
timestamp 1493745683
transform 1 0 332 0 1 450
box -3 -3 3 3
use $$M2_M1  $$M2_M1_119
timestamp 1493745683
transform 1 0 332 0 1 447
box -2 -2 2 2
use $$M3_M2  $$M3_M2_115
timestamp 1493745683
transform 1 0 316 0 1 440
box -3 -3 3 3
use $$M3_M2  $$M3_M2_117
timestamp 1493745683
transform 1 0 340 0 1 400
box -3 -3 3 3
use $$M2_M1  $$M2_M1_121
timestamp 1493745683
transform 1 0 396 0 1 400
box -2 -2 2 2
use $$M3_M2  $$M3_M2_118
timestamp 1493745683
transform 1 0 396 0 1 400
box -3 -3 3 3
use $$M2_M1  $$M2_M1_122
timestamp 1493745683
transform 1 0 404 0 1 400
box -2 -2 2 2
use $$M2_M1  $$M2_M1_120
timestamp 1493745683
transform 1 0 420 0 1 463
box -2 -2 2 2
use $$M3_M2  $$M3_M2_116
timestamp 1493745683
transform 1 0 428 0 1 410
box -3 -3 3 3
use $$M2_M1_1500_1500_3_1  $$M2_M1_1500_1500_3_1_10
timestamp 1493745683
transform 1 0 37 0 1 390
box -7 -2 7 2
use INVX2  INVX2_9
timestamp 1493745683
transform 1 0 80 0 -1 490
box -9 -3 26 105
use FILL  FILL_66
timestamp 1493745683
transform 1 0 96 0 -1 490
box -8 -3 16 105
use OAI21X1  OAI21X1_4
timestamp 1493745683
transform 1 0 104 0 -1 490
box -8 -3 34 105
use AOI21X1  AOI21X1_2
timestamp 1493745683
transform -1 0 168 0 -1 490
box -7 -3 39 105
use FILL  FILL_68
timestamp 1493745683
transform 1 0 168 0 -1 490
box -8 -3 16 105
use OAI21X1  OAI21X1_5
timestamp 1493745683
transform 1 0 176 0 -1 490
box -8 -3 34 105
use FILL  FILL_70
timestamp 1493745683
transform 1 0 208 0 -1 490
box -8 -3 16 105
use INVX1  INVX1_0
timestamp 1493147875
transform -1 0 232 0 -1 490
box -9 -3 26 105
use $$M3_M2  $$M3_M2_119
timestamp 1493745683
transform 1 0 244 0 1 390
box -3 -3 3 3
use NAND3X1  NAND3X1_3
timestamp 1493745683
transform 1 0 232 0 -1 490
box -8 -3 40 105
use FILL  FILL_80
timestamp 1493745683
transform 1 0 264 0 -1 490
box -8 -3 16 105
use FILL  FILL_81
timestamp 1493745683
transform 1 0 272 0 -1 490
box -8 -3 16 105
use FILL  FILL_82
timestamp 1493745683
transform 1 0 280 0 -1 490
box -8 -3 16 105
use FILL  FILL_83
timestamp 1493745683
transform 1 0 288 0 -1 490
box -8 -3 16 105
use $$M3_M2  $$M3_M2_139
timestamp 1493745683
transform 1 0 308 0 1 390
box -3 -3 3 3
use FILL  FILL_84
timestamp 1493745683
transform 1 0 296 0 -1 490
box -8 -3 16 105
use DFFPOSX1  DFFPOSX1_3
timestamp 1493147875
transform 1 0 304 0 -1 490
box -8 -3 104 105
use FILL  FILL_87
timestamp 1493745683
transform 1 0 400 0 -1 490
box -8 -3 16 105
use INVX1  INVX1_1
timestamp 1493147875
transform -1 0 424 0 -1 490
box -9 -3 26 105
use FILL  FILL_88
timestamp 1493745683
transform 1 0 424 0 -1 490
box -8 -3 16 105
use FILL  FILL_89
timestamp 1493745683
transform 1 0 432 0 -1 490
box -8 -3 16 105
use FILL  FILL_90
timestamp 1493745683
transform 1 0 440 0 -1 490
box -8 -3 16 105
use FILL  FILL_91
timestamp 1493745683
transform 1 0 448 0 -1 490
box -8 -3 16 105
use FILL  FILL_92
timestamp 1493745683
transform 1 0 456 0 -1 490
box -8 -3 16 105
use FILL  FILL_93
timestamp 1493745683
transform 1 0 464 0 -1 490
box -8 -3 16 105
use FILL  FILL_94
timestamp 1493745683
transform 1 0 472 0 -1 490
box -8 -3 16 105
use FILL  FILL_95
timestamp 1493745683
transform 1 0 480 0 -1 490
box -8 -3 16 105
use FILL  FILL_96
timestamp 1493745683
transform 1 0 488 0 -1 490
box -8 -3 16 105
use FILL  FILL_97
timestamp 1493745683
transform 1 0 496 0 -1 490
box -8 -3 16 105
use $$M2_M1_1500_1500_3_1  $$M2_M1_1500_1500_3_1_12
timestamp 1493745683
transform 1 0 546 0 1 390
box -7 -2 7 2
use $$M3_M2  $$M3_M2_121
timestamp 1493745683
transform 1 0 100 0 1 340
box -3 -3 3 3
use $$M2_M1  $$M2_M1_123
timestamp 1493745683
transform 1 0 100 0 1 333
box -2 -2 2 2
use $$M2_M1  $$M2_M1_125
timestamp 1493745683
transform 1 0 84 0 1 313
box -2 -2 2 2
use $$M3_M2  $$M3_M2_123
timestamp 1493745683
transform 1 0 84 0 1 310
box -3 -3 3 3
use $$M2_M1  $$M2_M1_129
timestamp 1493745683
transform 1 0 92 0 1 300
box -2 -2 2 2
use $$M3_M2  $$M3_M2_124
timestamp 1493745683
transform 1 0 108 0 1 310
box -3 -3 3 3
use $$M3_M2  $$M3_M2_120
timestamp 1493745683
transform 1 0 132 0 1 360
box -3 -3 3 3
use $$M3_M2  $$M3_M2_122
timestamp 1493745683
transform 1 0 124 0 1 340
box -3 -3 3 3
use $$M2_M1  $$M2_M1_124
timestamp 1493745683
transform 1 0 124 0 1 333
box -2 -2 2 2
use $$M3_M2  $$M3_M2_125
timestamp 1493745683
transform 1 0 156 0 1 350
box -3 -3 3 3
use $$M3_M2  $$M3_M2_126
timestamp 1493745683
transform 1 0 148 0 1 320
box -3 -3 3 3
use $$M2_M1  $$M2_M1_126
timestamp 1493745683
transform 1 0 156 0 1 321
box -2 -2 2 2
use $$M2_M1  $$M2_M1_127
timestamp 1493745683
transform 1 0 140 0 1 311
box -2 -2 2 2
use $$M2_M1  $$M2_M1_128
timestamp 1493745683
transform 1 0 148 0 1 310
box -2 -2 2 2
use $$M2_M1  $$M2_M1_130
timestamp 1493745683
transform 1 0 132 0 1 300
box -2 -2 2 2
use $$M3_M2  $$M3_M2_127
timestamp 1493745683
transform 1 0 132 0 1 300
box -3 -3 3 3
use $$M3_M2  $$M3_M2_128
timestamp 1493745683
transform 1 0 180 0 1 360
box -3 -3 3 3
use $$M3_M2  $$M3_M2_129
timestamp 1493745683
transform 1 0 172 0 1 340
box -3 -3 3 3
use $$M2_M1  $$M2_M1_131
timestamp 1493745683
transform 1 0 180 0 1 340
box -2 -2 2 2
use $$M3_M2  $$M3_M2_131
timestamp 1493745683
transform 1 0 172 0 1 320
box -3 -3 3 3
use $$M2_M1  $$M2_M1_133
timestamp 1493745683
transform 1 0 172 0 1 315
box -2 -2 2 2
use $$M3_M2  $$M3_M2_130
timestamp 1493745683
transform 1 0 188 0 1 340
box -3 -3 3 3
use $$M2_M1  $$M2_M1_132
timestamp 1493745683
transform 1 0 188 0 1 330
box -2 -2 2 2
use $$M3_M2  $$M3_M2_132
timestamp 1493745683
transform 1 0 204 0 1 360
box -3 -3 3 3
use $$M3_M2  $$M3_M2_133
timestamp 1493745683
transform 1 0 220 0 1 350
box -3 -3 3 3
use $$M2_M1  $$M2_M1_134
timestamp 1493745683
transform 1 0 228 0 1 350
box -2 -2 2 2
use $$M2_M1  $$M2_M1_135
timestamp 1493745683
transform 1 0 212 0 1 331
box -2 -2 2 2
use $$M2_M1  $$M2_M1_136
timestamp 1493745683
transform 1 0 220 0 1 330
box -2 -2 2 2
use $$M3_M2  $$M3_M2_134
timestamp 1493745683
transform 1 0 220 0 1 330
box -3 -3 3 3
use $$M3_M2  $$M3_M2_138
timestamp 1493745683
transform 1 0 236 0 1 350
box -3 -3 3 3
use $$M3_M2  $$M3_M2_135
timestamp 1493745683
transform 1 0 228 0 1 320
box -3 -3 3 3
use $$M3_M2  $$M3_M2_136
timestamp 1493745683
transform 1 0 212 0 1 300
box -3 -3 3 3
use $$M2_M1  $$M2_M1_137
timestamp 1493745683
transform 1 0 244 0 1 333
box -2 -2 2 2
use $$M2_M1  $$M2_M1_139
timestamp 1493745683
transform 1 0 236 0 1 320
box -2 -2 2 2
use $$M3_M2  $$M3_M2_137
timestamp 1493745683
transform 1 0 260 0 1 360
box -3 -3 3 3
use $$M2_M1  $$M2_M1_138
timestamp 1493745683
transform 1 0 260 0 1 328
box -2 -2 2 2
use $$M3_M2  $$M3_M2_140
timestamp 1493745683
transform 1 0 316 0 1 350
box -3 -3 3 3
use $$M2_M1  $$M2_M1_140
timestamp 1493745683
transform 1 0 292 0 1 331
box -2 -2 2 2
use $$M3_M2  $$M3_M2_141
timestamp 1493745683
transform 1 0 300 0 1 330
box -3 -3 3 3
use $$M2_M1  $$M2_M1_141
timestamp 1493745683
transform 1 0 308 0 1 331
box -2 -2 2 2
use $$M2_M1  $$M2_M1_142
timestamp 1493745683
transform 1 0 316 0 1 330
box -2 -2 2 2
use $$M3_M2  $$M3_M2_142
timestamp 1493745683
transform 1 0 276 0 1 320
box -3 -3 3 3
use $$M2_M1  $$M2_M1_143
timestamp 1493745683
transform 1 0 284 0 1 323
box -2 -2 2 2
use $$M3_M2  $$M3_M2_143
timestamp 1493745683
transform 1 0 292 0 1 320
box -3 -3 3 3
use $$M3_M2  $$M3_M2_144
timestamp 1493745683
transform 1 0 308 0 1 320
box -3 -3 3 3
use $$M2_M1  $$M2_M1_144
timestamp 1493745683
transform 1 0 260 0 1 311
box -2 -2 2 2
use $$M3_M2  $$M3_M2_148
timestamp 1493745683
transform 1 0 260 0 1 300
box -3 -3 3 3
use $$M2_M1  $$M2_M1_149
timestamp 1493745683
transform 1 0 308 0 1 310
box -2 -2 2 2
use $$M2_M1  $$M2_M1_150
timestamp 1493745683
transform 1 0 276 0 1 300
box -2 -2 2 2
use $$M2_M1  $$M2_M1_148
timestamp 1493745683
transform 1 0 324 0 1 312
box -2 -2 2 2
use $$M2_M1  $$M2_M1_145
timestamp 1493745683
transform 1 0 348 0 1 330
box -2 -2 2 2
use $$M3_M2  $$M3_M2_146
timestamp 1493745683
transform 1 0 340 0 1 320
box -3 -3 3 3
use $$M2_M1  $$M2_M1_151
timestamp 1493745683
transform 1 0 340 0 1 300
box -2 -2 2 2
use $$M3_M2  $$M3_M2_145
timestamp 1493745683
transform 1 0 364 0 1 340
box -3 -3 3 3
use $$M2_M1  $$M2_M1_146
timestamp 1493745683
transform 1 0 364 0 1 330
box -2 -2 2 2
use $$M3_M2  $$M3_M2_147
timestamp 1493745683
transform 1 0 356 0 1 320
box -3 -3 3 3
use $$M2_M1  $$M2_M1_153
timestamp 1493745683
transform 1 0 364 0 1 317
box -2 -2 2 2
use $$M2_M1  $$M2_M1_147
timestamp 1493745683
transform 1 0 372 0 1 330
box -2 -2 2 2
use $$M2_M1  $$M2_M1_152
timestamp 1493745683
transform 1 0 380 0 1 321
box -2 -2 2 2
use $$M3_M2  $$M3_M2_149
timestamp 1493745683
transform 1 0 404 0 1 350
box -3 -3 3 3
use $$M3_M2  $$M3_M2_150
timestamp 1493745683
transform 1 0 420 0 1 340
box -3 -3 3 3
use $$M3_M2  $$M3_M2_151
timestamp 1493745683
transform 1 0 412 0 1 330
box -3 -3 3 3
use $$M2_M1  $$M2_M1_154
timestamp 1493745683
transform 1 0 420 0 1 330
box -2 -2 2 2
use $$M2_M1  $$M2_M1_155
timestamp 1493745683
transform 1 0 404 0 1 320
box -2 -2 2 2
use $$M2_M1  $$M2_M1_156
timestamp 1493745683
transform 1 0 412 0 1 300
box -2 -2 2 2
use $$M3_M2  $$M3_M2_152
timestamp 1493745683
transform 1 0 420 0 1 300
box -3 -3 3 3
use $$M2_M1  $$M2_M1_157
timestamp 1493745683
transform 1 0 452 0 1 350
box -2 -2 2 2
use $$M2_M1  $$M2_M1_158
timestamp 1493745683
transform 1 0 436 0 1 340
box -2 -2 2 2
use $$M3_M2  $$M3_M2_153
timestamp 1493745683
transform 1 0 444 0 1 340
box -3 -3 3 3
use $$M2_M1  $$M2_M1_159
timestamp 1493745683
transform 1 0 444 0 1 334
box -2 -2 2 2
use $$M2_M1  $$M2_M1_160
timestamp 1493745683
transform 1 0 460 0 1 330
box -2 -2 2 2
use $$M3_M2  $$M3_M2_154
timestamp 1493745683
transform 1 0 460 0 1 330
box -3 -3 3 3
use $$M3_M2  $$M3_M2_155
timestamp 1493745683
transform 1 0 452 0 1 320
box -3 -3 3 3
use $$M3_M2  $$M3_M2_160
timestamp 1493745683
transform 1 0 484 0 1 330
box -3 -3 3 3
use $$M2_M1  $$M2_M1_161
timestamp 1493745683
transform 1 0 484 0 1 327
box -2 -2 2 2
use $$M2_M1  $$M2_M1_162
timestamp 1493745683
transform 1 0 492 0 1 300
box -2 -2 2 2
use $$M2_M1_1500_1500_3_1  $$M2_M1_1500_1500_3_1_11
timestamp 1493745683
transform 1 0 62 0 1 290
box -7 -2 7 2
use NOR2X1  NOR2X1_7
timestamp 1493745683
transform 1 0 80 0 1 290
box -8 -3 32 105
use FILL  FILL_98
timestamp 1493745683
transform -1 0 112 0 1 290
box -8 -3 16 105
use FILL  FILL_99
timestamp 1493745683
transform -1 0 120 0 1 290
box -8 -3 16 105
use NOR2X1  NOR2X1_8
timestamp 1493745683
transform -1 0 144 0 1 290
box -8 -3 32 105
use INVX2  INVX2_10
timestamp 1493745683
transform -1 0 160 0 1 290
box -9 -3 26 105
use FILL  FILL_103
timestamp 1493745683
transform -1 0 168 0 1 290
box -8 -3 16 105
use $$M3_M2  $$M3_M2_156
timestamp 1493745683
transform 1 0 196 0 1 290
box -3 -3 3 3
use NOR2X1  NOR2X1_9
timestamp 1493745683
transform 1 0 168 0 1 290
box -8 -3 32 105
use FILL  FILL_106
timestamp 1493745683
transform -1 0 200 0 1 290
box -8 -3 16 105
use OAI21X1  OAI21X1_6
timestamp 1493745683
transform 1 0 200 0 1 290
box -8 -3 34 105
use $$M3_M2  $$M3_M2_157
timestamp 1493745683
transform 1 0 244 0 1 290
box -3 -3 3 3
use FILL  FILL_108
timestamp 1493745683
transform -1 0 240 0 1 290
box -8 -3 16 105
use NOR2X1  NOR2X1_10
timestamp 1493745683
transform -1 0 264 0 1 290
box -8 -3 32 105
use INVX2  INVX2_11
timestamp 1493745683
transform 1 0 264 0 1 290
box -9 -3 26 105
use OAI22X1  OAI22X1_0
timestamp 1493745683
transform 1 0 280 0 1 290
box -8 -3 46 105
use FILL  FILL_110
timestamp 1493745683
transform -1 0 328 0 1 290
box -8 -3 16 105
use NOR2X1  NOR2X1_11
timestamp 1493745683
transform 1 0 328 0 1 290
box -8 -3 32 105
use FILL  FILL_115
timestamp 1493745683
transform -1 0 360 0 1 290
box -8 -3 16 105
use $$M3_M2  $$M3_M2_158
timestamp 1493745683
transform 1 0 380 0 1 290
box -3 -3 3 3
use INVX1  INVX1_2
timestamp 1493147875
transform 1 0 360 0 1 290
box -9 -3 26 105
use INVX2  INVX2_12
timestamp 1493745683
transform 1 0 376 0 1 290
box -9 -3 26 105
use FILL  FILL_118
timestamp 1493745683
transform -1 0 400 0 1 290
box -8 -3 16 105
use NOR2X1  NOR2X1_12
timestamp 1493745683
transform 1 0 400 0 1 290
box -8 -3 32 105
use $$M3_M2  $$M3_M2_159
timestamp 1493745683
transform 1 0 436 0 1 290
box -3 -3 3 3
use FILL  FILL_119
timestamp 1493745683
transform -1 0 432 0 1 290
box -8 -3 16 105
use NAND3X1  NAND3X1_4
timestamp 1493745683
transform 1 0 432 0 1 290
box -8 -3 40 105
use FILL  FILL_120
timestamp 1493745683
transform -1 0 472 0 1 290
box -8 -3 16 105
use FILL  FILL_121
timestamp 1493745683
transform -1 0 480 0 1 290
box -8 -3 16 105
use INVX2  INVX2_13
timestamp 1493745683
transform 1 0 480 0 1 290
box -9 -3 26 105
use FILL  FILL_122
timestamp 1493745683
transform -1 0 504 0 1 290
box -8 -3 16 105
use $$M2_M1_1500_1500_3_1  $$M2_M1_1500_1500_3_1_13
timestamp 1493745683
transform 1 0 521 0 1 290
box -7 -2 7 2
use $$M3_M2  $$M3_M2_161
timestamp 1493745683
transform 1 0 92 0 1 270
box -3 -3 3 3
use $$M2_M1  $$M2_M1_163
timestamp 1493745683
transform 1 0 92 0 1 263
box -2 -2 2 2
use $$M3_M2  $$M3_M2_162
timestamp 1493745683
transform 1 0 92 0 1 260
box -3 -3 3 3
use $$M3_M2  $$M3_M2_163
timestamp 1493745683
transform 1 0 108 0 1 260
box -3 -3 3 3
use $$M3_M2  $$M3_M2_164
timestamp 1493745683
transform 1 0 108 0 1 250
box -3 -3 3 3
use $$M2_M1  $$M2_M1_164
timestamp 1493745683
transform 1 0 108 0 1 247
box -2 -2 2 2
use $$M3_M2  $$M3_M2_165
timestamp 1493745683
transform 1 0 84 0 1 240
box -3 -3 3 3
use $$M2_M1  $$M2_M1_165
timestamp 1493745683
transform 1 0 100 0 1 240
box -2 -2 2 2
use $$M3_M2  $$M3_M2_166
timestamp 1493745683
transform 1 0 100 0 1 240
box -3 -3 3 3
use $$M3_M2  $$M3_M2_167
timestamp 1493745683
transform 1 0 84 0 1 200
box -3 -3 3 3
use $$M2_M1  $$M2_M1_166
timestamp 1493745683
transform 1 0 124 0 1 261
box -2 -2 2 2
use $$M3_M2  $$M3_M2_169
timestamp 1493745683
transform 1 0 124 0 1 250
box -3 -3 3 3
use $$M3_M2  $$M3_M2_168
timestamp 1493745683
transform 1 0 140 0 1 270
box -3 -3 3 3
use $$M3_M2  $$M3_M2_172
timestamp 1493745683
transform 1 0 156 0 1 270
box -3 -3 3 3
use $$M2_M1  $$M2_M1_167
timestamp 1493745683
transform 1 0 132 0 1 234
box -2 -2 2 2
use $$M3_M2  $$M3_M2_170
timestamp 1493745683
transform 1 0 132 0 1 230
box -3 -3 3 3
use $$M3_M2  $$M3_M2_171
timestamp 1493745683
transform 1 0 132 0 1 200
box -3 -3 3 3
use $$M2_M1  $$M2_M1_168
timestamp 1493745683
transform 1 0 164 0 1 253
box -2 -2 2 2
use $$M2_M1  $$M2_M1_169
timestamp 1493745683
transform 1 0 156 0 1 240
box -2 -2 2 2
use $$M3_M2  $$M3_M2_173
timestamp 1493745683
transform 1 0 164 0 1 240
box -3 -3 3 3
use $$M3_M2  $$M3_M2_174
timestamp 1493745683
transform 1 0 172 0 1 230
box -3 -3 3 3
use $$M2_M1  $$M2_M1_170
timestamp 1493745683
transform 1 0 212 0 1 248
box -2 -2 2 2
use $$M2_M1  $$M2_M1_171
timestamp 1493745683
transform 1 0 244 0 1 280
box -2 -2 2 2
use $$M2_M1  $$M2_M1_172
timestamp 1493745683
transform 1 0 236 0 1 255
box -2 -2 2 2
use $$M2_M1  $$M2_M1_173
timestamp 1493745683
transform 1 0 228 0 1 250
box -2 -2 2 2
use $$M3_M2  $$M3_M2_175
timestamp 1493745683
transform 1 0 228 0 1 250
box -3 -3 3 3
use $$M2_M1  $$M2_M1_174
timestamp 1493745683
transform 1 0 220 0 1 240
box -2 -2 2 2
use $$M3_M2  $$M3_M2_176
timestamp 1493745683
transform 1 0 220 0 1 240
box -3 -3 3 3
use $$M2_M1  $$M2_M1_175
timestamp 1493745683
transform 1 0 196 0 1 230
box -2 -2 2 2
use $$M3_M2  $$M3_M2_177
timestamp 1493745683
transform 1 0 212 0 1 230
box -3 -3 3 3
use $$M3_M2  $$M3_M2_178
timestamp 1493745683
transform 1 0 196 0 1 220
box -3 -3 3 3
use $$M2_M1  $$M2_M1_176
timestamp 1493745683
transform 1 0 188 0 1 200
box -2 -2 2 2
use $$M3_M2  $$M3_M2_179
timestamp 1493745683
transform 1 0 188 0 1 200
box -3 -3 3 3
use $$M3_M2  $$M3_M2_180
timestamp 1493745683
transform 1 0 236 0 1 220
box -3 -3 3 3
use $$M3_M2  $$M3_M2_181
timestamp 1493745683
transform 1 0 252 0 1 270
box -3 -3 3 3
use $$M2_M1  $$M2_M1_178
timestamp 1493745683
transform 1 0 268 0 1 250
box -2 -2 2 2
use $$M3_M2  $$M3_M2_186
timestamp 1493745683
transform 1 0 260 0 1 240
box -3 -3 3 3
use $$M2_M1  $$M2_M1_182
timestamp 1493745683
transform 1 0 252 0 1 230
box -2 -2 2 2
use $$M3_M2  $$M3_M2_182
timestamp 1493745683
transform 1 0 284 0 1 270
box -3 -3 3 3
use $$M2_M1  $$M2_M1_177
timestamp 1493745683
transform 1 0 300 0 1 280
box -2 -2 2 2
use $$M3_M2  $$M3_M2_187
timestamp 1493745683
transform 1 0 292 0 1 240
box -3 -3 3 3
use $$M2_M1  $$M2_M1_183
timestamp 1493745683
transform 1 0 292 0 1 230
box -2 -2 2 2
use $$M3_M2  $$M3_M2_183
timestamp 1493745683
transform 1 0 324 0 1 270
box -3 -3 3 3
use $$M2_M1  $$M2_M1_179
timestamp 1493745683
transform 1 0 324 0 1 253
box -2 -2 2 2
use $$M3_M2  $$M3_M2_184
timestamp 1493745683
transform 1 0 340 0 1 270
box -3 -3 3 3
use $$M3_M2  $$M3_M2_185
timestamp 1493745683
transform 1 0 356 0 1 270
box -3 -3 3 3
use $$M2_M1  $$M2_M1_181
timestamp 1493745683
transform 1 0 332 0 1 240
box -2 -2 2 2
use $$M2_M1  $$M2_M1_180
timestamp 1493745683
transform 1 0 340 0 1 243
box -2 -2 2 2
use $$M3_M2  $$M3_M2_188
timestamp 1493745683
transform 1 0 324 0 1 230
box -3 -3 3 3
use $$M2_M1  $$M2_M1_184
timestamp 1493745683
transform 1 0 348 0 1 230
box -2 -2 2 2
use $$M3_M2  $$M3_M2_189
timestamp 1493745683
transform 1 0 348 0 1 230
box -3 -3 3 3
use $$M2_M1  $$M2_M1_185
timestamp 1493745683
transform 1 0 356 0 1 200
box -2 -2 2 2
use $$M3_M2  $$M3_M2_190
timestamp 1493745683
transform 1 0 380 0 1 270
box -3 -3 3 3
use $$M3_M2  $$M3_M2_191
timestamp 1493745683
transform 1 0 372 0 1 250
box -3 -3 3 3
use $$M2_M1  $$M2_M1_186
timestamp 1493745683
transform 1 0 380 0 1 250
box -2 -2 2 2
use $$M2_M1  $$M2_M1_187
timestamp 1493745683
transform 1 0 372 0 1 200
box -2 -2 2 2
use $$M3_M2  $$M3_M2_193
timestamp 1493745683
transform 1 0 396 0 1 260
box -3 -3 3 3
use $$M3_M2  $$M3_M2_195
timestamp 1493745683
transform 1 0 396 0 1 250
box -3 -3 3 3
use $$M2_M1  $$M2_M1_189
timestamp 1493745683
transform 1 0 396 0 1 241
box -2 -2 2 2
use $$M2_M1  $$M2_M1_188
timestamp 1493745683
transform 1 0 420 0 1 260
box -2 -2 2 2
use $$M3_M2  $$M3_M2_194
timestamp 1493745683
transform 1 0 420 0 1 260
box -3 -3 3 3
use $$M3_M2  $$M3_M2_196
timestamp 1493745683
transform 1 0 412 0 1 230
box -3 -3 3 3
use $$M2_M1  $$M2_M1_191
timestamp 1493745683
transform 1 0 420 0 1 230
box -2 -2 2 2
use $$M2_M1  $$M2_M1_192
timestamp 1493745683
transform 1 0 404 0 1 200
box -2 -2 2 2
use $$M3_M2  $$M3_M2_192
timestamp 1493745683
transform 1 0 444 0 1 270
box -3 -3 3 3
use $$M2_M1  $$M2_M1_190
timestamp 1493745683
transform 1 0 444 0 1 255
box -2 -2 2 2
use $$M2_M1  $$M2_M1_193
timestamp 1493745683
transform 1 0 436 0 1 200
box -2 -2 2 2
use $$M3_M2  $$M3_M2_197
timestamp 1493745683
transform 1 0 436 0 1 200
box -3 -3 3 3
use $$M2_M1_1500_1500_3_1  $$M2_M1_1500_1500_3_1_14
timestamp 1493745683
transform 1 0 37 0 1 190
box -7 -2 7 2
use FILL  FILL_100
timestamp 1493745683
transform 1 0 80 0 -1 290
box -8 -3 16 105
use NOR2X1  NOR2X1_13
timestamp 1493745683
transform 1 0 88 0 -1 290
box -8 -3 32 105
use FILL  FILL_101
timestamp 1493745683
transform 1 0 112 0 -1 290
box -8 -3 16 105
use NOR2X1  NOR2X1_14
timestamp 1493745683
transform 1 0 120 0 -1 290
box -8 -3 32 105
use FILL  FILL_102
timestamp 1493745683
transform 1 0 144 0 -1 290
box -8 -3 16 105
use INVX2  INVX2_14
timestamp 1493745683
transform -1 0 168 0 -1 290
box -9 -3 26 105
use FILL  FILL_104
timestamp 1493745683
transform 1 0 168 0 -1 290
box -8 -3 16 105
use FILL  FILL_105
timestamp 1493745683
transform 1 0 176 0 -1 290
box -8 -3 16 105
use NAND3X1  NAND3X1_5
timestamp 1493745683
transform -1 0 216 0 -1 290
box -8 -3 40 105
use FILL  FILL_107
timestamp 1493745683
transform 1 0 216 0 -1 290
box -8 -3 16 105
use $$M3_M2  $$M3_M2_198
timestamp 1493745683
transform 1 0 244 0 1 190
box -3 -3 3 3
use INVX2  INVX2_15
timestamp 1493745683
transform -1 0 240 0 -1 290
box -9 -3 26 105
use FILL  FILL_109
timestamp 1493745683
transform 1 0 240 0 -1 290
box -8 -3 16 105
use $$M3_M2  $$M3_M2_199
timestamp 1493745683
transform 1 0 268 0 1 190
box -3 -3 3 3
use NAND2X1  NAND2X1_1
timestamp 1493745683
transform -1 0 272 0 -1 290
box -8 -3 32 105
use FILL  FILL_111
timestamp 1493745683
transform 1 0 272 0 -1 290
box -8 -3 16 105
use FILL  FILL_112
timestamp 1493745683
transform 1 0 280 0 -1 290
box -8 -3 16 105
use NAND2X1  NAND2X1_2
timestamp 1493745683
transform -1 0 312 0 -1 290
box -8 -3 32 105
use FILL  FILL_113
timestamp 1493745683
transform 1 0 312 0 -1 290
box -8 -3 16 105
use FILL  FILL_114
timestamp 1493745683
transform 1 0 320 0 -1 290
box -8 -3 16 105
use NAND3X1  NAND3X1_6
timestamp 1493745683
transform 1 0 328 0 -1 290
box -8 -3 40 105
use FILL  FILL_116
timestamp 1493745683
transform 1 0 360 0 -1 290
box -8 -3 16 105
use INVX2  INVX2_16
timestamp 1493745683
transform -1 0 384 0 -1 290
box -9 -3 26 105
use FILL  FILL_117
timestamp 1493745683
transform 1 0 384 0 -1 290
box -8 -3 16 105
use NOR2X1  NOR2X1_15
timestamp 1493745683
transform -1 0 416 0 -1 290
box -8 -3 32 105
use FILL  FILL_123
timestamp 1493745683
transform 1 0 416 0 -1 290
box -8 -3 16 105
use $$M3_M2  $$M3_M2_200
timestamp 1493745683
transform 1 0 452 0 1 190
box -3 -3 3 3
use NAND2X1  NAND2X1_3
timestamp 1493745683
transform -1 0 448 0 -1 290
box -8 -3 32 105
use FILL  FILL_124
timestamp 1493745683
transform 1 0 448 0 -1 290
box -8 -3 16 105
use FILL  FILL_125
timestamp 1493745683
transform 1 0 456 0 -1 290
box -8 -3 16 105
use FILL  FILL_126
timestamp 1493745683
transform 1 0 464 0 -1 290
box -8 -3 16 105
use FILL  FILL_127
timestamp 1493745683
transform 1 0 472 0 -1 290
box -8 -3 16 105
use FILL  FILL_128
timestamp 1493745683
transform 1 0 480 0 -1 290
box -8 -3 16 105
use FILL  FILL_129
timestamp 1493745683
transform 1 0 488 0 -1 290
box -8 -3 16 105
use FILL  FILL_130
timestamp 1493745683
transform 1 0 496 0 -1 290
box -8 -3 16 105
use $$M2_M1_1500_1500_3_1  $$M2_M1_1500_1500_3_1_15
timestamp 1493745683
transform 1 0 546 0 1 190
box -7 -2 7 2
use $$M2_M1_1500_1500_3_1  $$M2_M1_1500_1500_3_1_16
timestamp 1493745683
transform 1 0 62 0 1 90
box -7 -2 7 2
use $$M2_M1  $$M2_M1_194
timestamp 1493745683
transform 1 0 92 0 1 170
box -2 -2 2 2
use $$M3_M2  $$M3_M2_201
timestamp 1493745683
transform 1 0 92 0 1 170
box -3 -3 3 3
use FILL  FILL_131
timestamp 1493745683
transform -1 0 88 0 1 90
box -8 -3 16 105
use $$M2_M1  $$M2_M1_195
timestamp 1493745683
transform 1 0 100 0 1 121
box -2 -2 2 2
use $$M3_M2  $$M3_M2_202
timestamp 1493745683
transform 1 0 100 0 1 120
box -3 -3 3 3
use $$M2_M1  $$M2_M1_196
timestamp 1493745683
transform 1 0 108 0 1 100
box -2 -2 2 2
use INVX2  INVX2_17
timestamp 1493745683
transform -1 0 104 0 1 90
box -9 -3 26 105
use $$M3_M2  $$M3_M2_204
timestamp 1493745683
transform 1 0 124 0 1 150
box -3 -3 3 3
use $$M2_M1  $$M2_M1_199
timestamp 1493745683
transform 1 0 124 0 1 127
box -2 -2 2 2
use $$M3_M2  $$M3_M2_203
timestamp 1493745683
transform 1 0 148 0 1 170
box -3 -3 3 3
use $$M2_M1  $$M2_M1_197
timestamp 1493745683
transform 1 0 148 0 1 150
box -2 -2 2 2
use $$M3_M2  $$M3_M2_205
timestamp 1493745683
transform 1 0 148 0 1 150
box -3 -3 3 3
use $$M2_M1  $$M2_M1_198
timestamp 1493745683
transform 1 0 140 0 1 130
box -2 -2 2 2
use $$M3_M2  $$M3_M2_206
timestamp 1493745683
transform 1 0 140 0 1 130
box -3 -3 3 3
use INVX2  INVX2_18
timestamp 1493745683
transform -1 0 120 0 1 90
box -9 -3 26 105
use $$M2_M1  $$M2_M1_200
timestamp 1493745683
transform 1 0 132 0 1 125
box -2 -2 2 2
use $$M3_M2  $$M3_M2_207
timestamp 1493745683
transform 1 0 132 0 1 120
box -3 -3 3 3
use FILL  FILL_132
timestamp 1493745683
transform -1 0 128 0 1 90
box -8 -3 16 105
use NAND2X1  NAND2X1_4
timestamp 1493745683
transform 1 0 128 0 1 90
box -8 -3 32 105
use $$M3_M2  $$M3_M2_208
timestamp 1493745683
transform 1 0 196 0 1 170
box -3 -3 3 3
use $$M3_M2  $$M3_M2_209
timestamp 1493745683
transform 1 0 180 0 1 160
box -3 -3 3 3
use $$M2_M1  $$M2_M1_201
timestamp 1493745683
transform 1 0 164 0 1 150
box -2 -2 2 2
use $$M3_M2  $$M3_M2_210
timestamp 1493745683
transform 1 0 164 0 1 150
box -3 -3 3 3
use $$M2_M1  $$M2_M1_202
timestamp 1493745683
transform 1 0 172 0 1 150
box -2 -2 2 2
use FILL  FILL_133
timestamp 1493745683
transform -1 0 160 0 1 90
box -8 -3 16 105
use $$M2_M1  $$M2_M1_203
timestamp 1493745683
transform 1 0 180 0 1 140
box -2 -2 2 2
use $$M3_M2  $$M3_M2_214
timestamp 1493745683
transform 1 0 172 0 1 130
box -3 -3 3 3
use $$M3_M2  $$M3_M2_216
timestamp 1493745683
transform 1 0 172 0 1 110
box -3 -3 3 3
use $$M2_M1  $$M2_M1_207
timestamp 1493745683
transform 1 0 196 0 1 130
box -2 -2 2 2
use NAND3X1  NAND3X1_7
timestamp 1493745683
transform -1 0 192 0 1 90
box -8 -3 40 105
use FILL  FILL_134
timestamp 1493745683
transform -1 0 200 0 1 90
box -8 -3 16 105
use $$M2_M1  $$M2_M1_204
timestamp 1493745683
transform 1 0 260 0 1 180
box -2 -2 2 2
use $$M3_M2  $$M3_M2_211
timestamp 1493745683
transform 1 0 252 0 1 170
box -3 -3 3 3
use $$M3_M2  $$M3_M2_212
timestamp 1493745683
transform 1 0 244 0 1 160
box -3 -3 3 3
use $$M3_M2  $$M3_M2_213
timestamp 1493745683
transform 1 0 236 0 1 150
box -3 -3 3 3
use $$M2_M1  $$M2_M1_205
timestamp 1493745683
transform 1 0 212 0 1 138
box -2 -2 2 2
use $$M2_M1  $$M2_M1_206
timestamp 1493745683
transform 1 0 228 0 1 135
box -2 -2 2 2
use $$M3_M2  $$M3_M2_215
timestamp 1493745683
transform 1 0 228 0 1 130
box -3 -3 3 3
use $$M2_M1  $$M2_M1_208
timestamp 1493745683
transform 1 0 236 0 1 127
box -2 -2 2 2
use $$M2_M1  $$M2_M1_209
timestamp 1493745683
transform 1 0 212 0 1 110
box -2 -2 2 2
use $$M3_M2  $$M3_M2_217
timestamp 1493745683
transform 1 0 212 0 1 110
box -3 -3 3 3
use $$M3_M2  $$M3_M2_218
timestamp 1493745683
transform 1 0 236 0 1 110
box -3 -3 3 3
use OAI22X1  OAI22X1_1
timestamp 1493745683
transform -1 0 240 0 1 90
box -8 -3 46 105
use $$M2_M1  $$M2_M1_211
timestamp 1493745683
transform 1 0 252 0 1 119
box -2 -2 2 2
use FILL  FILL_135
timestamp 1493745683
transform -1 0 248 0 1 90
box -8 -3 16 105
use $$M2_M1  $$M2_M1_210
timestamp 1493745683
transform 1 0 268 0 1 130
box -2 -2 2 2
use $$M3_M2  $$M3_M2_219
timestamp 1493745683
transform 1 0 268 0 1 130
box -3 -3 3 3
use NOR2X1  NOR2X1_16
timestamp 1493745683
transform 1 0 248 0 1 90
box -8 -3 32 105
use $$M3_M2  $$M3_M2_220
timestamp 1493745683
transform 1 0 300 0 1 170
box -3 -3 3 3
use $$M2_M1  $$M2_M1_212
timestamp 1493745683
transform 1 0 287 0 1 160
box -2 -2 2 2
use $$M3_M2  $$M3_M2_221
timestamp 1493745683
transform 1 0 287 0 1 160
box -3 -3 3 3
use $$M3_M2  $$M3_M2_222
timestamp 1493745683
transform 1 0 284 0 1 140
box -3 -3 3 3
use $$M2_M1  $$M2_M1_213
timestamp 1493745683
transform 1 0 284 0 1 136
box -2 -2 2 2
use FILL  FILL_136
timestamp 1493745683
transform -1 0 280 0 1 90
box -8 -3 16 105
use $$M2_M1  $$M2_M1_214
timestamp 1493745683
transform 1 0 300 0 1 117
box -2 -2 2 2
use $$M3_M2  $$M3_M2_224
timestamp 1493745683
transform 1 0 316 0 1 140
box -3 -3 3 3
use $$M2_M1  $$M2_M1_215
timestamp 1493745683
transform 1 0 340 0 1 150
box -2 -2 2 2
use $$M3_M2  $$M3_M2_223
timestamp 1493745683
transform 1 0 340 0 1 150
box -3 -3 3 3
use $$M2_M1  $$M2_M1_217
timestamp 1493745683
transform 1 0 316 0 1 127
box -2 -2 2 2
use $$M2_M1  $$M2_M1_216
timestamp 1493745683
transform 1 0 324 0 1 133
box -2 -2 2 2
use $$M3_M2  $$M3_M2_225
timestamp 1493745683
transform 1 0 324 0 1 130
box -3 -3 3 3
use $$M3_M2  $$M3_M2_227
timestamp 1493745683
transform 1 0 308 0 1 110
box -3 -3 3 3
use NOR2X1  NOR2X1_17
timestamp 1493745683
transform -1 0 304 0 1 90
box -8 -3 32 105
use FILL  FILL_137
timestamp 1493745683
transform -1 0 312 0 1 90
box -8 -3 16 105
use $$M3_M2  $$M3_M2_228
timestamp 1493745683
transform 1 0 332 0 1 100
box -3 -3 3 3
use $$M3_M2  $$M3_M2_226
timestamp 1493745683
transform 1 0 348 0 1 130
box -3 -3 3 3
use $$M2_M1  $$M2_M1_218
timestamp 1493745683
transform 1 0 340 0 1 100
box -2 -2 2 2
use $$M3_M2  $$M3_M2_229
timestamp 1493745683
transform 1 0 340 0 1 90
box -3 -3 3 3
use OAI21X1  OAI21X1_7
timestamp 1493745683
transform 1 0 312 0 1 90
box -8 -3 34 105
use $$M2_M1  $$M2_M1_220
timestamp 1493745683
transform 1 0 356 0 1 127
box -2 -2 2 2
use FILL  FILL_138
timestamp 1493745683
transform -1 0 352 0 1 90
box -8 -3 16 105
use FILL  FILL_139
timestamp 1493745683
transform -1 0 360 0 1 90
box -8 -3 16 105
use $$M3_M2  $$M3_M2_230
timestamp 1493745683
transform 1 0 388 0 1 170
box -3 -3 3 3
use $$M2_M1  $$M2_M1_219
timestamp 1493745683
transform 1 0 380 0 1 150
box -2 -2 2 2
use $$M3_M2  $$M3_M2_231
timestamp 1493745683
transform 1 0 380 0 1 150
box -3 -3 3 3
use $$M2_M1  $$M2_M1_222
timestamp 1493745683
transform 1 0 412 0 1 137
box -2 -2 2 2
use $$M2_M1  $$M2_M1_223
timestamp 1493745683
transform 1 0 404 0 1 123
box -2 -2 2 2
use $$M2_M1  $$M2_M1_224
timestamp 1493745683
transform 1 0 388 0 1 111
box -2 -2 2 2
use $$M2_M1  $$M2_M1_221
timestamp 1493745683
transform 1 0 372 0 1 100
box -2 -2 2 2
use $$M3_M2  $$M3_M2_232
timestamp 1493745683
transform 1 0 372 0 1 100
box -3 -3 3 3
use $$M3_M2  $$M3_M2_233
timestamp 1493745683
transform 1 0 388 0 1 100
box -3 -3 3 3
use $$M3_M2  $$M3_M2_234
timestamp 1493745683
transform 1 0 372 0 1 90
box -3 -3 3 3
use INVX2  INVX2_19
timestamp 1493745683
transform 1 0 360 0 1 90
box -9 -3 26 105
use FILL  FILL_140
timestamp 1493745683
transform -1 0 384 0 1 90
box -8 -3 16 105
use AOI21X1  AOI21X1_3
timestamp 1493745683
transform -1 0 416 0 1 90
box -7 -3 39 105
use FILL  FILL_141
timestamp 1493745683
transform -1 0 424 0 1 90
box -8 -3 16 105
use FILL  FILL_142
timestamp 1493745683
transform -1 0 432 0 1 90
box -8 -3 16 105
use FILL  FILL_143
timestamp 1493745683
transform -1 0 440 0 1 90
box -8 -3 16 105
use $$M2_M1  $$M2_M1_225
timestamp 1493745683
transform 1 0 452 0 1 127
box -2 -2 2 2
use FILL  FILL_144
timestamp 1493745683
transform -1 0 448 0 1 90
box -8 -3 16 105
use $$M2_M1  $$M2_M1_226
timestamp 1493745683
transform 1 0 460 0 1 100
box -2 -2 2 2
use INVX2  INVX2_20
timestamp 1493745683
transform 1 0 448 0 1 90
box -9 -3 26 105
use FILL  FILL_145
timestamp 1493745683
transform -1 0 472 0 1 90
box -8 -3 16 105
use FILL  FILL_146
timestamp 1493745683
transform -1 0 480 0 1 90
box -8 -3 16 105
use FILL  FILL_147
timestamp 1493745683
transform -1 0 488 0 1 90
box -8 -3 16 105
use FILL  FILL_148
timestamp 1493745683
transform -1 0 496 0 1 90
box -8 -3 16 105
use FILL  FILL_149
timestamp 1493745683
transform -1 0 504 0 1 90
box -8 -3 16 105
use $$M2_M1_1500_1500_3_1  $$M2_M1_1500_1500_3_1_17
timestamp 1493745683
transform 1 0 521 0 1 90
box -7 -2 7 2
use $$M2_M1_1500_1500_3_3  $$M2_M1_1500_1500_3_3_4
timestamp 1493745683
transform 1 0 62 0 1 72
box -7 -7 7 7
use $$M3_M2  $$M3_M2_235
timestamp 1493745683
transform 1 0 116 0 1 80
box -3 -3 3 3
use $$M2_M1_1500_1500_3_3  $$M2_M1_1500_1500_3_3_5
timestamp 1493745683
transform 1 0 521 0 1 72
box -7 -7 7 7
use $$M3_M2  $$M3_M2_236
timestamp 1493745683
transform 1 0 108 0 1 60
box -3 -3 3 3
use $$M3_M2  $$M3_M2_237
timestamp 1493745683
transform 1 0 460 0 1 60
box -3 -3 3 3
use $$M2_M1_1500_1500_3_3  $$M2_M1_1500_1500_3_3_6
timestamp 1493745683
transform 1 0 37 0 1 47
box -7 -7 7 7
use $$M2_M1_1500_1500_3_3  $$M2_M1_1500_1500_3_3_7
timestamp 1493745683
transform 1 0 546 0 1 47
box -7 -7 7 7
use $$M2_M1  $$M2_M1_227
timestamp 1493745683
transform 1 0 268 0 1 30
box -2 -2 2 2
use $$M2_M1  $$M2_M1_228
timestamp 1493745683
transform 1 0 500 0 1 30
box -2 -2 2 2
<< labels >>
flabel metal3 2 80 2 80 4 FreeSans 26 0 0 0 reset
flabel metal3 2 200 2 200 4 FreeSans 26 0 0 0 irwrite[3]
flabel metal3 2 920 2 920 4 FreeSans 26 0 0 0 clk
flabel metal3 2 300 2 300 4 FreeSans 26 0 0 0 irwrite[0]
flabel metal3 2 330 2 330 4 FreeSans 26 0 0 0 iord
flabel metal3 2 270 2 270 4 FreeSans 26 0 0 0 irwrite[1]
flabel metal3 2 230 2 230 4 FreeSans 26 0 0 0 irwrite[2]
flabel metal3 2 130 2 130 4 FreeSans 26 0 0 0 regwrite
flabel metal3 2 170 2 170 4 FreeSans 26 0 0 0 regdst
flabel metal3 2 60 2 60 4 FreeSans 26 0 0 0 memtoreg
flabel metal2 132 978 132 978 4 FreeSans 26 0 0 0 op[2]
flabel metal2 44 978 44 978 4 FreeSans 26 0 0 0 op[5]
flabel metal2 100 978 100 978 4 FreeSans 26 0 0 0 op[3]
flabel metal2 68 978 68 978 4 FreeSans 26 0 0 0 op[4]
flabel metal2 172 978 172 978 4 FreeSans 26 0 0 0 op[1]
flabel metal2 204 978 204 978 4 FreeSans 26 0 0 0 op[0]
flabel metal2 332 978 332 978 4 FreeSans 26 0 0 0 memwrite
flabel metal3 581 920 581 920 4 FreeSans 26 0 0 0 aluop[0]
flabel metal3 581 60 581 60 4 FreeSans 26 0 0 0 aluop[1]
flabel metal2 268 1 268 1 4 FreeSans 26 0 0 0 pcsrc[0]
flabel metal2 204 1 204 1 4 FreeSans 26 0 0 0 alusrcb[1]
flabel metal2 332 1 332 1 4 FreeSans 26 0 0 0 pcsrc[1]
flabel metal2 172 1 172 1 4 FreeSans 26 0 0 0 alusrcb[0]
flabel metal2 236 1 236 1 4 FreeSans 26 0 0 0 alusrca
flabel metal2 404 1 404 1 4 FreeSans 26 0 0 0 zero
flabel metal2 372 1 372 1 4 FreeSans 26 0 0 0 pcen
rlabel metal1 374 930 374 930 1 Vdd!
rlabel metal1 374 905 374 905 1 Gnd!
<< end >>
