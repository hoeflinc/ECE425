magic
tech scmos
timestamp 1493754735
<< m2contact >>
rect 1295 2494 1299 2498
rect 273 1340 277 1344
<< metal2 >>
rect 487 2552 491 2556
rect 241 1344 245 1845
rect 904 1541 908 1815
rect 924 1719 928 2512
rect 934 1749 938 2530
rect 944 1789 948 2521
rect 966 2439 970 2594
rect 1006 2494 1010 2539
rect 1030 2497 1034 2548
rect 1062 2497 1066 2557
rect 1095 2494 1099 2566
rect 1134 2497 1138 2575
rect 1166 2497 1170 2584
rect 1631 1720 1635 2421
rect 1653 1737 1657 2405
rect 1678 1756 1682 2389
rect 1705 1775 1709 2378
rect 1752 1794 1756 2354
rect 1787 1833 1791 2339
rect 1819 1813 1823 2326
rect 1884 1911 1888 2435
rect 2019 2329 2023 2339
rect 2090 2328 2094 2354
rect 2154 2320 2158 2378
rect 2218 2329 2222 2389
rect 2290 2326 2294 2405
rect 2354 2322 2358 2421
rect 250 1380 254 1537
rect 265 1343 269 1523
rect 922 1446 926 1573
rect 305 1344 309 1376
rect 942 1354 946 1685
rect 950 1344 954 1645
rect 958 1527 962 1595
rect 1914 1579 1918 1947
rect 966 1424 970 1575
rect 1135 1460 1138 1518
rect 1167 1470 1170 1519
rect 1199 1480 1202 1519
rect 1231 1490 1234 1517
rect 1295 1500 1298 1518
rect 1335 1510 1338 1519
rect 1321 1344 1325 1456
rect 1353 1342 1357 1466
rect 1529 1340 1533 1476
rect 1681 1344 1685 1486
rect 1713 1344 1717 1496
rect 1769 1344 1773 1506
rect 1937 1343 1941 1516
rect 1962 1364 1966 1854
rect 2019 1849 2020 1855
rect 1992 1676 1996 1716
rect 1992 1341 1996 1672
rect 2000 1692 2004 1733
rect 2000 1339 2004 1688
rect 2019 1374 2023 1849
rect 2032 1340 2036 1752
rect 2048 1340 2052 1771
rect 2065 1340 2069 1790
rect 2090 1384 2094 1853
rect 2154 1394 2158 1852
rect 2184 1340 2188 1809
rect 2218 1404 2222 1856
rect 2291 1855 2294 1861
rect 2250 1344 2254 1829
rect 2290 1414 2294 1855
rect 2529 1672 2533 1688
rect 2528 1346 2532 1442
rect 2224 1340 2254 1344
rect 1391 1067 1395 1124
rect 2077 1036 2081 1064
rect 2640 1015 2644 1032
<< m3contact >>
rect 287 2769 291 2773
rect 383 2594 387 2598
rect 966 2594 970 2598
rect 471 2584 475 2588
rect 463 2575 467 2579
rect 455 2566 459 2570
rect 447 2557 451 2561
rect 439 2548 443 2552
rect 431 2539 435 2543
rect 487 2530 491 2534
rect 934 2530 938 2534
rect 671 2521 675 2525
rect 303 2512 307 2516
rect 924 2512 928 2516
rect 241 1845 245 1849
rect 904 1815 908 1819
rect 944 2521 948 2525
rect 1166 2584 1170 2588
rect 1134 2575 1138 2579
rect 1095 2566 1099 2570
rect 1062 2557 1066 2561
rect 1030 2548 1034 2552
rect 1006 2539 1010 2543
rect 966 2435 970 2439
rect 1884 2435 1888 2439
rect 944 1785 948 1789
rect 1631 2421 1635 2425
rect 934 1745 938 1749
rect 924 1715 928 1719
rect 1653 2405 1657 2409
rect 1678 2389 1682 2393
rect 1705 2378 1709 2382
rect 1752 2354 1756 2358
rect 1787 2339 1791 2343
rect 1787 1829 1791 1833
rect 1819 2326 1823 2330
rect 2354 2421 2358 2425
rect 2290 2405 2294 2409
rect 2218 2389 2222 2393
rect 2154 2378 2158 2382
rect 2090 2354 2094 2358
rect 2019 2339 2023 2343
rect 1966 2326 1970 2330
rect 1884 1907 1888 1911
rect 1914 1947 1918 1951
rect 1819 1809 1823 1813
rect 1752 1790 1756 1794
rect 1705 1771 1709 1775
rect 1678 1752 1682 1756
rect 1653 1733 1657 1737
rect 1631 1716 1635 1720
rect 942 1685 946 1689
rect 250 1537 254 1541
rect 904 1537 908 1541
rect 922 1573 926 1577
rect 250 1376 254 1380
rect 265 1523 269 1527
rect 922 1442 926 1446
rect 305 1376 309 1380
rect 942 1350 946 1354
rect 950 1645 954 1649
rect 958 1595 962 1599
rect 958 1523 962 1527
rect 966 1575 970 1579
rect 1914 1575 1918 1579
rect 1366 1516 1370 1520
rect 1937 1516 1941 1520
rect 1335 1506 1339 1510
rect 1769 1506 1773 1510
rect 1295 1496 1299 1500
rect 1713 1496 1717 1500
rect 1231 1486 1235 1490
rect 1681 1486 1685 1490
rect 1199 1476 1203 1480
rect 1529 1476 1533 1480
rect 1167 1466 1171 1470
rect 1353 1466 1357 1470
rect 1135 1456 1139 1460
rect 1321 1456 1325 1460
rect 966 1420 970 1424
rect 950 1340 954 1344
rect 2000 1733 2004 1737
rect 1962 1360 1966 1364
rect 1992 1716 1996 1720
rect 1992 1672 1996 1676
rect 2000 1688 2004 1692
rect 2065 1790 2069 1794
rect 2048 1771 2052 1775
rect 2019 1370 2023 1374
rect 2032 1752 2036 1756
rect 2154 1390 2158 1394
rect 2184 1809 2188 1813
rect 2090 1380 2094 1384
rect 2218 1400 2222 1404
rect 2250 1829 2254 1833
rect 2529 1688 2533 1692
rect 2472 1672 2476 1676
rect 2290 1410 2294 1414
rect 2528 1442 2532 1446
rect 1391 1124 1395 1128
rect 2592 1124 2596 1128
rect 1409 1064 1413 1068
rect 2077 1064 2081 1068
rect 2077 1032 2081 1036
rect 2640 1032 2644 1036
<< metal3 >>
rect 382 2598 971 2599
rect 382 2594 383 2598
rect 387 2594 966 2598
rect 970 2594 971 2598
rect 382 2593 971 2594
rect 470 2588 1171 2589
rect 470 2584 471 2588
rect 475 2584 1166 2588
rect 1170 2584 1171 2588
rect 470 2583 1171 2584
rect 462 2579 1139 2580
rect 462 2575 463 2579
rect 467 2575 1134 2579
rect 1138 2575 1139 2579
rect 462 2574 1139 2575
rect 454 2570 1100 2571
rect 454 2566 455 2570
rect 459 2566 1095 2570
rect 1099 2566 1100 2570
rect 454 2565 1100 2566
rect 446 2561 1067 2562
rect 446 2557 447 2561
rect 451 2557 1062 2561
rect 1066 2557 1067 2561
rect 446 2556 1067 2557
rect 438 2552 1035 2553
rect 438 2548 439 2552
rect 443 2548 1030 2552
rect 1034 2548 1035 2552
rect 438 2547 1035 2548
rect 430 2543 1011 2544
rect 430 2539 431 2543
rect 435 2539 1006 2543
rect 1010 2539 1011 2543
rect 430 2538 1011 2539
rect 486 2534 939 2535
rect 486 2530 487 2534
rect 491 2530 934 2534
rect 938 2530 939 2534
rect 486 2529 939 2530
rect 670 2525 949 2526
rect 670 2521 671 2525
rect 675 2521 944 2525
rect 948 2521 949 2525
rect 670 2520 949 2521
rect 302 2516 929 2517
rect 302 2512 303 2516
rect 307 2512 924 2516
rect 928 2512 929 2516
rect 302 2511 929 2512
rect 965 2439 971 2440
rect 965 2435 966 2439
rect 970 2435 971 2439
rect 965 2434 971 2435
rect 1549 2439 1889 2440
rect 1549 2435 1884 2439
rect 1888 2435 1889 2439
rect 1549 2434 1889 2435
rect 1630 2425 2359 2426
rect 1630 2421 1631 2425
rect 1635 2421 2354 2425
rect 2358 2421 2359 2425
rect 1630 2420 2359 2421
rect 1652 2409 2295 2410
rect 1652 2405 1653 2409
rect 1657 2405 2290 2409
rect 2294 2405 2295 2409
rect 1652 2404 2295 2405
rect 1677 2393 2223 2394
rect 1677 2389 1678 2393
rect 1682 2389 2218 2393
rect 2222 2389 2223 2393
rect 1677 2388 2223 2389
rect 1704 2382 2159 2383
rect 1704 2378 1705 2382
rect 1709 2378 2154 2382
rect 2158 2378 2159 2382
rect 1704 2377 2159 2378
rect 1751 2358 2095 2359
rect 1751 2354 1752 2358
rect 1756 2354 2090 2358
rect 2094 2354 2095 2358
rect 1751 2353 2095 2354
rect 1786 2343 2024 2344
rect 1786 2339 1787 2343
rect 1791 2339 2019 2343
rect 2023 2339 2024 2343
rect 1786 2338 2024 2339
rect 1818 2330 1971 2331
rect 1818 2326 1819 2330
rect 1823 2326 1966 2330
rect 1970 2326 1971 2330
rect 1818 2325 1971 2326
rect 1913 1951 1921 1952
rect 1913 1947 1914 1951
rect 1918 1947 1921 1951
rect 1913 1946 1921 1947
rect 1883 1911 1921 1912
rect 1883 1907 1884 1911
rect 1888 1907 1921 1911
rect 1883 1906 1921 1907
rect 240 1849 965 1850
rect 240 1845 241 1849
rect 245 1845 965 1849
rect 240 1844 965 1845
rect 1786 1833 2255 1834
rect 1786 1829 1787 1833
rect 1791 1829 2250 1833
rect 2254 1829 2255 1833
rect 1786 1828 2255 1829
rect 903 1819 965 1820
rect 903 1815 904 1819
rect 908 1815 965 1819
rect 903 1814 965 1815
rect 1818 1813 2189 1814
rect 1818 1809 1819 1813
rect 1823 1809 2184 1813
rect 2188 1809 2189 1813
rect 1818 1808 2189 1809
rect 1751 1794 2070 1795
rect 1751 1790 1752 1794
rect 1756 1790 2065 1794
rect 2069 1790 2070 1794
rect 943 1789 965 1790
rect 1751 1789 2070 1790
rect 943 1785 944 1789
rect 948 1785 965 1789
rect 943 1784 965 1785
rect 1704 1775 2053 1776
rect 1704 1771 1705 1775
rect 1709 1771 2048 1775
rect 2052 1771 2053 1775
rect 1704 1770 2053 1771
rect 1677 1756 2037 1757
rect 1677 1752 1678 1756
rect 1682 1752 2032 1756
rect 2036 1752 2037 1756
rect 1677 1751 2037 1752
rect 933 1749 966 1750
rect 933 1745 934 1749
rect 938 1745 966 1749
rect 933 1744 966 1745
rect 1652 1737 2005 1738
rect 1652 1733 1653 1737
rect 1657 1733 2000 1737
rect 2004 1733 2005 1737
rect 1652 1732 2005 1733
rect 1630 1720 1997 1721
rect 923 1719 965 1720
rect 923 1715 924 1719
rect 928 1715 965 1719
rect 1630 1716 1631 1720
rect 1635 1716 1992 1720
rect 1996 1716 1997 1720
rect 1630 1715 1997 1716
rect 923 1714 965 1715
rect 1999 1692 2534 1693
rect 941 1689 965 1690
rect 941 1685 942 1689
rect 946 1685 965 1689
rect 1999 1688 2000 1692
rect 2004 1688 2529 1692
rect 2533 1688 2534 1692
rect 1999 1687 2534 1688
rect 941 1684 965 1685
rect 1991 1676 2477 1677
rect 1991 1672 1992 1676
rect 1996 1672 2472 1676
rect 2476 1672 2477 1676
rect 1991 1671 2477 1672
rect 949 1649 965 1650
rect 949 1645 950 1649
rect 954 1645 965 1649
rect 949 1644 965 1645
rect 957 1599 965 1600
rect 957 1595 958 1599
rect 962 1595 965 1599
rect 957 1594 965 1595
rect 965 1579 971 1580
rect 965 1575 966 1579
rect 970 1575 971 1579
rect 965 1574 971 1575
rect 1549 1579 1919 1580
rect 1549 1575 1914 1579
rect 1918 1575 1919 1579
rect 1549 1574 1919 1575
rect 249 1541 909 1542
rect 249 1537 250 1541
rect 254 1537 904 1541
rect 908 1537 909 1541
rect 249 1536 909 1537
rect 264 1527 963 1528
rect 264 1523 265 1527
rect 269 1523 958 1527
rect 962 1523 963 1527
rect 264 1522 963 1523
rect 1365 1520 1942 1521
rect 1365 1516 1366 1520
rect 1370 1516 1937 1520
rect 1941 1516 1942 1520
rect 1365 1515 1942 1516
rect 1334 1510 1774 1511
rect 1334 1506 1335 1510
rect 1339 1506 1769 1510
rect 1773 1506 1774 1510
rect 1334 1505 1774 1506
rect 1294 1500 1718 1501
rect 1294 1496 1295 1500
rect 1299 1496 1713 1500
rect 1717 1496 1718 1500
rect 1294 1495 1718 1496
rect 1230 1490 1686 1491
rect 1230 1486 1231 1490
rect 1235 1486 1681 1490
rect 1685 1486 1686 1490
rect 1230 1485 1686 1486
rect 1198 1480 1534 1481
rect 1198 1476 1199 1480
rect 1203 1476 1529 1480
rect 1533 1476 1534 1480
rect 1198 1475 1534 1476
rect 1166 1470 1358 1471
rect 1166 1466 1167 1470
rect 1171 1466 1353 1470
rect 1357 1466 1358 1470
rect 1166 1465 1358 1466
rect 1134 1460 1326 1461
rect 1134 1456 1135 1460
rect 1139 1456 1321 1460
rect 1325 1456 1326 1460
rect 1134 1455 1326 1456
rect 921 1446 2533 1447
rect 921 1442 922 1446
rect 926 1442 2528 1446
rect 2532 1442 2533 1446
rect 921 1441 2533 1442
rect 507 1424 971 1425
rect 507 1420 966 1424
rect 970 1420 971 1424
rect 507 1419 971 1420
rect 517 1414 2295 1415
rect 517 1410 2290 1414
rect 2294 1410 2295 1414
rect 517 1409 2295 1410
rect 522 1404 2223 1405
rect 522 1400 2218 1404
rect 2222 1400 2223 1404
rect 522 1399 2223 1400
rect 538 1394 2159 1395
rect 538 1390 2154 1394
rect 2158 1390 2159 1394
rect 538 1389 2159 1390
rect 547 1384 2095 1385
rect 249 1380 310 1381
rect 249 1376 250 1380
rect 254 1376 305 1380
rect 309 1376 310 1380
rect 547 1380 2090 1384
rect 2094 1380 2095 1384
rect 547 1379 2095 1380
rect 249 1375 310 1376
rect 551 1374 2024 1375
rect 551 1370 2019 1374
rect 2023 1370 2024 1374
rect 551 1369 2024 1370
rect 675 1364 1967 1365
rect 675 1360 1962 1364
rect 1966 1360 1967 1364
rect 675 1359 1967 1360
rect 708 1354 947 1355
rect 708 1350 942 1354
rect 946 1350 947 1354
rect 708 1349 947 1350
rect 712 1344 955 1345
rect 712 1340 950 1344
rect 954 1340 955 1344
rect 712 1339 955 1340
rect 1390 1128 2597 1129
rect 1390 1124 1391 1128
rect 1395 1124 2592 1128
rect 2596 1124 2597 1128
rect 1390 1123 2597 1124
rect 1408 1068 2082 1069
rect 1408 1064 1409 1068
rect 1413 1064 2077 1068
rect 2081 1064 2082 1068
rect 1408 1063 2082 1064
rect 2076 1036 2645 1037
rect 2076 1032 2077 1036
rect 2081 1032 2640 1036
rect 2644 1032 2645 1036
rect 2076 1031 2645 1032
rect 233 880 237 884
rect 233 870 237 874
rect 233 860 237 864
rect 230 770 234 774
rect 230 760 234 764
rect 230 750 234 754
rect 230 660 234 664
rect 230 650 234 654
rect 230 640 234 644
rect 230 550 234 554
rect 230 540 234 544
rect 230 530 234 534
rect 230 440 234 444
rect 230 430 234 434
rect 230 420 234 424
rect 230 330 234 334
rect 230 320 234 324
rect 230 310 234 314
rect 230 220 234 224
rect 230 210 234 214
rect 230 200 234 204
rect 230 110 234 114
rect 230 100 234 104
rect 230 90 234 94
use mips_fsm  mips_fsm_0
timestamp 1493746172
transform 1 0 965 0 1 1517
box 0 0 584 980
use aludec  aludec_0
timestamp 1493749612
transform 1 0 1921 0 1 1849
box 0 0 850 480
use datapath_new  datapath_new_0
timestamp 1493661823
transform 1 0 -279 0 1 32
box 279 -32 3123 2811
<< labels >>
rlabel metal3 233 880 237 884 1 memdata7
rlabel metal3 233 870 237 874 1 writedata7
rlabel metal3 233 860 237 864 1 adr7
rlabel metal3 230 770 234 774 1 memdata6
rlabel metal3 230 760 234 764 1 writedata6
rlabel metal3 230 750 234 754 1 adr6
rlabel metal3 230 660 234 664 1 memdata5
rlabel metal3 230 650 234 654 1 writedata5
rlabel metal3 230 640 234 644 1 adr5
rlabel metal3 230 550 234 554 1 memdata4
rlabel metal3 230 540 234 544 1 writedata4
rlabel metal3 230 530 234 534 1 adr4
rlabel metal3 230 440 234 444 1 memdata3
rlabel metal3 230 430 234 434 1 writedata3
rlabel metal3 230 420 234 424 1 adr3
rlabel metal3 230 330 234 334 1 memdata2
rlabel metal3 230 320 234 324 1 writedata2
rlabel metal3 230 310 234 314 1 adr2
rlabel metal3 230 220 234 224 1 memdata1
rlabel metal3 230 200 234 204 1 adr1
rlabel metal3 230 110 234 114 1 memdata0
rlabel metal3 230 100 234 104 1 writedata0
rlabel metal3 230 90 234 94 1 adr0
rlabel metal3 230 210 234 214 1 writedata1
rlabel m2contact 273 1340 277 1344 1 ph2
rlabel metal3 957 1594 965 1600 1 reset
rlabel m2contact 1295 2494 1299 2498 1 memwrite
rlabel m3contact 287 2769 291 2773 1 ph1
rlabel metal3 1575 2437 1575 2437 1 aluop0
rlabel metal3 1603 1577 1603 1577 1 aluop1
rlabel metal3 1246 1469 1247 1469 1 alusrcb1
rlabel metal3 1257 1458 1257 1458 1 alusrcb0
rlabel metal3 1499 1497 1499 1497 1 pcsrc1
rlabel metal3 1154 2586 1154 2586 1 op0
rlabel metal3 1127 2577 1127 2577 1 op1
rlabel metal3 1089 2569 1089 2569 1 op2
rlabel metal3 1057 2559 1057 2559 1 op3
rlabel metal3 1025 2550 1025 2550 1 op4
rlabel metal3 1001 2542 1001 2542 1 op5
rlabel metal3 959 1817 959 1817 1 irwrite0
rlabel metal3 960 1787 960 1787 1 irwrite1
rlabel metal3 959 1747 959 1747 1 irwrite2
rlabel metal3 958 1717 958 1717 1 irwrite3
<< end >>
