magic
tech scmos
timestamp 1488310061
<< m2contact >>
rect -7 -7 7 7
<< end >>
