magic
tech scmos
timestamp 1493147875
<< m2contact >>
rect -7 -7 7 7
<< end >>
