magic
tech scmos
timestamp 1485891256
<< nwell >>
rect -12 -4 32 23
<< ntransistor >>
rect -1 -38 1 -26
rect 10 -38 12 -26
rect 18 -38 20 -26
<< ptransistor >>
rect -1 2 1 10
rect 10 2 12 10
rect 18 2 20 10
<< ndiffusion >>
rect -2 -38 -1 -26
rect 1 -38 10 -26
rect 12 -38 18 -26
rect 20 -38 21 -26
<< pdiffusion >>
rect -2 2 -1 10
rect 1 2 5 10
rect 9 2 10 10
rect 12 2 13 10
rect 17 2 18 10
rect 20 2 21 10
<< ndcontact >>
rect -6 -38 -2 -26
rect 21 -38 25 -26
<< pdcontact >>
rect -6 2 -2 10
rect 5 2 9 10
rect 13 2 17 10
rect 21 2 25 10
<< psubstratepcontact >>
rect 29 -46 33 -42
<< nsubstratencontact >>
rect 22 14 26 18
<< polysilicon >>
rect -1 10 1 12
rect 10 10 12 12
rect 18 10 20 12
rect -1 -2 1 2
rect -1 -26 1 -6
rect 10 -10 12 2
rect 10 -26 12 -14
rect 18 -18 20 2
rect 18 -26 20 -22
rect -1 -40 1 -38
rect 10 -40 12 -38
rect 18 -40 20 -38
<< polycontact >>
rect -3 -6 1 -2
rect 8 -14 12 -10
rect 16 -22 20 -18
<< metal1 >>
rect -17 14 22 18
rect 26 14 36 18
rect -6 10 -2 14
rect 13 10 17 14
rect 5 -2 9 2
rect 21 -2 25 2
rect -17 -6 -3 -2
rect 5 -6 28 -2
rect -17 -14 8 -10
rect 24 -13 28 -6
rect 24 -17 36 -13
rect -17 -22 16 -18
rect 24 -26 28 -17
rect 25 -30 28 -26
rect -6 -42 -2 -38
rect -17 -46 29 -42
rect 33 -46 36 -42
<< labels >>
rlabel metal1 -17 -6 -17 -6 3 A
rlabel metal1 -17 -14 -17 -14 3 B
rlabel metal1 -17 -22 -17 -22 3 C
rlabel metal1 -6 14 -6 14 4 Vdd!
rlabel metal1 34 -15 34 -15 7 Y
rlabel metal1 -17 -42 -17 -42 2 Gnd!
<< end >>
