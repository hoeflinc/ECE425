magic
tech scmos
timestamp 1488306862
<< m2contact >>
rect -7 -7 7 7
<< end >>
