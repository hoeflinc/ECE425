magic
tech scmos
timestamp 1493063752
<< metal1 >>
rect 276 970 284 978
<< m2contact >>
rect 253 799 257 803
rect 326 772 330 776
rect 326 662 330 666
rect 326 552 330 556
rect 326 442 330 446
rect -17 367 -13 371
rect 326 332 330 336
rect 326 222 330 226
rect 326 112 330 116
<< metal2 >>
rect 246 922 250 986
rect -25 676 -21 711
rect -9 690 -5 782
rect -25 536 -21 562
rect -25 456 -21 491
rect -9 470 -5 532
rect -25 236 -21 271
rect -9 250 -5 342
rect -25 16 -21 51
rect -9 30 -5 122
rect 54 38 58 888
rect 62 38 66 888
rect 94 53 98 888
rect 110 37 114 888
rect 127 55 131 888
rect 254 877 258 926
rect 286 922 290 986
rect 254 872 258 873
rect 158 719 162 825
rect 253 767 257 799
rect 158 609 162 715
rect 158 499 162 605
rect 158 389 162 495
rect 158 279 162 385
rect 158 169 162 275
rect 158 59 162 165
rect 270 46 274 873
rect 278 834 282 922
rect 294 877 298 926
rect 302 53 306 922
rect 318 38 322 873
rect 326 776 330 826
rect 326 666 330 716
rect 326 556 330 606
rect 326 446 330 496
rect 326 336 330 386
rect 326 226 330 276
rect 326 116 330 166
rect 335 56 339 763
rect 350 60 354 830
<< m3contact >>
rect -9 782 -5 786
rect -25 672 -21 676
rect -25 562 -21 566
rect -25 532 -21 536
rect -9 532 -5 536
rect -25 452 -21 456
rect -9 342 -5 346
rect -25 232 -21 236
rect -9 122 -5 126
rect 270 922 274 926
rect 278 922 282 926
rect 254 873 258 877
rect 270 873 274 877
rect 253 763 257 767
rect 127 51 131 55
rect 158 51 162 55
rect 294 873 298 877
rect 302 922 306 926
rect 310 922 314 926
rect 278 830 282 834
rect 318 873 322 877
rect 350 830 354 834
rect 335 763 339 767
rect 326 52 330 56
rect 335 52 339 56
rect -25 12 -21 16
<< metal3 >>
rect 269 926 283 927
rect 269 922 270 926
rect 274 922 278 926
rect 282 922 283 926
rect 269 921 283 922
rect 301 926 315 927
rect 301 922 302 926
rect 306 922 310 926
rect 314 922 315 926
rect 301 921 315 922
rect 253 877 275 878
rect 253 873 254 877
rect 258 873 270 877
rect 274 873 275 877
rect 253 872 275 873
rect 293 877 323 878
rect 293 873 294 877
rect 298 873 318 877
rect 322 873 323 877
rect 293 872 323 873
rect -31 851 -5 857
rect -31 841 -5 847
rect 277 834 355 835
rect 277 830 278 834
rect 282 830 350 834
rect 354 830 355 834
rect 277 829 355 830
rect -31 786 -5 787
rect -31 782 -9 786
rect -31 781 -5 782
rect 252 767 340 768
rect 252 763 253 767
rect 257 763 335 767
rect 339 763 340 767
rect 252 762 340 763
rect -31 741 -5 747
rect -31 731 -5 737
rect -31 676 -5 677
rect -31 672 -25 676
rect -21 672 -5 676
rect -31 671 -5 672
rect -31 631 -5 637
rect -31 621 -5 627
rect -31 566 -5 567
rect -31 562 -25 566
rect -21 562 -5 566
rect -31 561 -5 562
rect -26 536 -4 537
rect -26 532 -25 536
rect -21 532 -9 536
rect -5 532 -4 536
rect -26 531 -4 532
rect -31 521 -5 527
rect -31 511 -5 517
rect -31 456 -5 457
rect -31 452 -25 456
rect -21 452 -5 456
rect -31 451 -5 452
rect -31 411 -5 417
rect -31 401 -5 407
rect -31 346 -5 347
rect -31 342 -9 346
rect -31 341 -5 342
rect -31 301 -5 307
rect -31 291 -5 297
rect -31 236 -5 237
rect -31 232 -25 236
rect -21 232 -5 236
rect -31 231 -5 232
rect -31 191 -5 197
rect -31 181 -5 187
rect -31 126 -5 127
rect -31 122 -9 126
rect -31 121 -5 122
rect -31 81 -5 87
rect -31 71 -5 77
rect 325 56 340 57
rect 126 55 163 56
rect 126 51 127 55
rect 131 51 158 55
rect 162 51 163 55
rect 325 52 326 56
rect 330 52 335 56
rect 339 52 340 56
rect 325 51 340 52
rect 126 50 163 51
rect -31 16 -5 17
rect -31 12 -25 16
rect -21 12 -5 16
rect -31 11 -5 12
use invbuf_4x  invbuf_4x_0
timestamp 1484532969
transform 1 0 246 0 1 884
box -6 -4 34 96
use invbuf_4x  invbuf_4x_1
timestamp 1484532969
transform 1 0 286 0 1 884
box -6 -4 34 96
use yzdetect_8  yzdetect_8_0
timestamp 1484534894
transform 1 0 -25 0 1 4
box -8 -4 28 756
use alt_alu_slice  alt_alu_slice_0
array 0 0 55 0 7 110
timestamp 1492981790
transform 1 0 0 0 1 0
box -5 0 377 100
<< labels >>
rlabel metal2 129 886 129 886 5 op2
rlabel metal2 56 886 56 886 5 op6
rlabel metal2 64 886 64 886 5 op5
rlabel metal2 96 886 96 886 5 op4
rlabel metal2 112 886 112 886 5 op3
rlabel metal2 248 984 248 984 5 op0
rlabel metal2 288 984 288 984 5 op1
rlabel metal3 -28 84 -28 84 3 a_0_
rlabel metal3 -29 74 -29 74 3 b_0_
rlabel metal3 -29 14 -29 14 3 result_0_
rlabel metal3 -29 194 -29 194 3 a_1_
rlabel metal3 -29 184 -29 184 3 b_1_
rlabel metal3 -29 124 -29 124 3 result_1_
rlabel metal3 -29 304 -29 304 3 a_2_
rlabel metal3 -29 294 -29 294 3 b_2_
rlabel metal3 -29 234 -29 234 3 result_2_
rlabel metal3 -29 414 -29 414 3 a_3_
rlabel metal3 -29 404 -29 404 3 b_3_
rlabel metal3 -28 344 -28 344 3 result_3_
rlabel metal3 -28 524 -28 524 3 a_4_
rlabel metal3 -28 514 -28 514 3 b_4_
rlabel metal3 -27 454 -27 454 1 result_4_
rlabel metal3 -29 634 -29 634 3 a_5_
rlabel metal3 -29 624 -29 624 3 b_5_
rlabel metal3 -28 564 -28 564 3 result_5_
rlabel metal3 -29 744 -29 744 3 a_6_
rlabel metal3 -29 734 -29 734 3 b_6_
rlabel metal3 -29 674 -29 674 3 result_6_
rlabel metal3 -29 854 -29 854 3 a_7_
rlabel metal3 -29 844 -29 844 3 b_7_
rlabel metal3 -29 784 -29 784 3 result_7_
rlabel m2contact -17 367 -13 371 1 zero
<< end >>
