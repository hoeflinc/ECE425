magic
tech scmos
timestamp 1493661823
<< metal1 >>
rect 576 2465 1096 2473
rect 576 2375 1096 2383
rect 576 2355 1096 2363
rect 703 2311 710 2315
rect 887 2311 894 2315
rect 576 2265 1096 2273
rect 576 2245 1096 2253
rect 703 2201 718 2205
rect 887 2201 902 2205
rect 576 2155 1096 2163
rect 576 2135 1096 2143
rect 703 2091 726 2095
rect 887 2091 910 2095
rect 1071 2091 1078 2095
rect 576 2045 1096 2053
rect 576 2025 1096 2033
rect 703 1981 734 1985
rect 1071 1981 1086 1985
rect 576 1935 1096 1943
rect 576 1915 1096 1923
rect 703 1871 742 1875
rect 1071 1871 1094 1875
rect 576 1825 1096 1833
rect 576 1805 1096 1813
rect 703 1761 750 1765
rect 887 1761 918 1765
rect 576 1715 1096 1723
rect 576 1695 1096 1703
rect 887 1651 926 1655
rect 576 1605 1096 1613
rect 576 1585 1096 1593
rect 887 1541 934 1545
rect 576 1495 1096 1503
rect 279 1302 3033 1304
rect 343 1298 2969 1302
rect 279 1296 3033 1298
rect 817 1248 827 1252
rect 369 1212 3123 1214
rect 433 1208 3059 1212
rect 369 1206 3123 1208
rect 820 1198 856 1202
rect 876 1198 888 1202
rect 279 1192 3033 1194
rect 343 1188 2969 1192
rect 279 1186 3033 1188
rect 369 1102 3123 1104
rect 433 1098 3059 1102
rect 369 1096 3123 1098
rect 820 1088 872 1092
rect 279 1082 3033 1084
rect 343 1078 2969 1082
rect 279 1076 3033 1078
rect 369 992 3123 994
rect 433 988 3059 992
rect 369 986 3123 988
rect 279 972 3033 974
rect 343 968 2969 972
rect 279 966 3033 968
rect 369 882 3123 884
rect 433 878 3059 882
rect 369 876 3123 878
rect 279 862 2231 864
rect 343 858 2231 862
rect 279 856 2231 858
rect 2479 862 3033 864
rect 2479 858 2969 862
rect 2479 856 3033 858
rect 856 816 875 820
rect 856 813 860 816
rect 1808 815 1812 819
rect 1801 811 1812 815
rect 2032 812 2067 816
rect 2032 808 2036 812
rect 369 772 2231 774
rect 433 771 2231 772
rect 433 768 1624 771
rect 369 767 1624 768
rect 1628 767 2231 771
rect 369 766 2231 767
rect 2479 772 3123 774
rect 2479 768 3059 772
rect 2479 766 3123 768
rect 1668 757 1672 761
rect 279 752 2199 754
rect 343 748 2199 752
rect 279 746 2199 748
rect 2479 752 3033 754
rect 2479 748 2969 752
rect 2479 746 3033 748
rect 856 706 875 710
rect 856 703 860 706
rect 1808 705 1812 709
rect 1801 701 1812 705
rect 2032 702 2067 706
rect 2032 698 2036 702
rect 1660 693 1664 697
rect 369 662 2199 664
rect 433 661 2199 662
rect 433 658 1624 661
rect 369 657 1624 658
rect 1628 657 2199 661
rect 369 656 2199 657
rect 2479 662 3123 664
rect 2479 658 3059 662
rect 2479 656 3123 658
rect 1668 647 1672 651
rect 279 642 2199 644
rect 343 638 2199 642
rect 279 636 2199 638
rect 2479 642 3033 644
rect 2479 638 2969 642
rect 2479 636 3033 638
rect 856 596 875 600
rect 705 592 712 596
rect 856 593 860 596
rect 1808 595 1812 599
rect 1801 591 1812 595
rect 2032 592 2067 596
rect 2032 588 2036 592
rect 1660 583 1664 587
rect 369 552 2199 554
rect 433 551 2199 552
rect 433 548 1624 551
rect 369 547 1624 548
rect 1628 547 2199 551
rect 369 546 2199 547
rect 2479 552 3123 554
rect 2479 548 3059 552
rect 2479 546 3123 548
rect 1668 537 1672 541
rect 279 532 2199 534
rect 343 528 2199 532
rect 279 526 2199 528
rect 2479 532 3033 534
rect 2479 528 2969 532
rect 2479 526 3033 528
rect 856 486 875 490
rect 705 482 720 486
rect 856 483 860 486
rect 1808 485 1812 489
rect 1801 481 1812 485
rect 2032 482 2067 486
rect 2032 478 2036 482
rect 1660 473 1664 477
rect 369 442 2199 444
rect 433 441 2199 442
rect 433 438 1624 441
rect 369 437 1624 438
rect 1628 437 2199 441
rect 369 436 2199 437
rect 2479 442 3123 444
rect 2479 438 3059 442
rect 2479 436 3123 438
rect 1668 427 1672 431
rect 279 422 2199 424
rect 343 418 2199 422
rect 279 416 2199 418
rect 2479 422 3033 424
rect 2479 418 2969 422
rect 2479 416 3033 418
rect 856 376 875 380
rect 705 372 728 376
rect 856 373 860 376
rect 1808 375 1812 379
rect 1801 371 1812 375
rect 2032 372 2067 376
rect 2032 368 2036 372
rect 1660 363 1664 367
rect 2201 363 2216 367
rect 369 333 581 334
rect 758 333 2199 334
rect 369 332 2199 333
rect 433 331 2199 332
rect 433 328 1624 331
rect 369 327 1624 328
rect 1628 327 2199 331
rect 369 326 2199 327
rect 2479 332 3123 334
rect 2479 328 3059 332
rect 2479 326 3123 328
rect 573 325 925 326
rect 1668 317 1672 321
rect 279 312 2199 314
rect 343 308 2199 312
rect 279 306 2199 308
rect 2479 312 3033 314
rect 2479 308 2969 312
rect 2479 306 3033 308
rect 856 266 875 270
rect 705 262 736 266
rect 856 263 860 266
rect 1808 265 1812 269
rect 1801 261 1812 265
rect 2032 262 2067 266
rect 2032 258 2036 262
rect 1660 253 1664 257
rect 369 222 2199 224
rect 433 221 2199 222
rect 433 218 1624 221
rect 369 217 1624 218
rect 1628 217 2199 221
rect 369 216 2199 217
rect 2479 222 3123 224
rect 2479 218 3059 222
rect 2479 216 3123 218
rect 1668 207 1672 211
rect 279 202 2199 204
rect 343 198 2199 202
rect 279 196 2199 198
rect 2479 202 3033 204
rect 2479 198 2969 202
rect 2479 196 3033 198
rect 856 156 875 160
rect 704 152 744 156
rect 856 153 860 156
rect 1808 155 1812 159
rect 1801 151 1812 155
rect 2032 152 2067 156
rect 2032 148 2036 152
rect 369 112 2199 114
rect 433 111 2199 112
rect 433 108 1624 111
rect 369 107 1624 108
rect 1628 107 1672 111
rect 1676 107 2199 111
rect 369 106 2199 107
rect 2479 112 3123 114
rect 2479 108 3059 112
rect 2479 106 3123 108
rect 279 92 2199 94
rect 343 91 2199 92
rect 343 88 1624 91
rect 279 87 1624 88
rect 1628 87 2199 91
rect 279 86 2199 87
rect 2479 92 3033 94
rect 2479 88 2969 92
rect 2479 86 3033 88
rect 856 46 875 50
rect 704 42 752 46
rect 856 43 860 46
rect 1808 45 1812 49
rect 1801 41 1812 45
rect 2032 42 2067 46
rect 2032 38 2036 42
rect 1660 33 1664 37
rect 369 2 2199 4
rect 433 1 2199 2
rect 433 -2 1672 1
rect 369 -3 1672 -2
rect 1676 -3 2199 1
rect 369 -4 2199 -3
rect 2479 2 3123 4
rect 2479 -2 3059 2
rect 2479 -4 3123 -2
<< m2contact >>
rect 710 2311 714 2315
rect 894 2311 898 2315
rect 718 2201 722 2205
rect 902 2201 906 2205
rect 726 2091 730 2095
rect 910 2091 914 2095
rect 1078 2091 1082 2095
rect 734 1981 738 1985
rect 1086 1981 1090 1985
rect 742 1871 746 1875
rect 1094 1871 1098 1875
rect 750 1761 754 1765
rect 918 1761 922 1765
rect 926 1651 930 1655
rect 2751 1640 2755 1644
rect 2808 1640 2812 1644
rect 934 1541 938 1545
rect 279 1298 343 1302
rect 2969 1298 3033 1302
rect 369 1208 433 1212
rect 3059 1208 3123 1212
rect 816 1198 820 1202
rect 856 1198 860 1202
rect 872 1198 876 1202
rect 888 1198 892 1202
rect 279 1188 343 1192
rect 2969 1188 3033 1192
rect 369 1098 433 1102
rect 3059 1098 3123 1102
rect 816 1088 820 1092
rect 872 1088 876 1092
rect 279 1078 343 1082
rect 2969 1078 3033 1082
rect 369 988 433 992
rect 3059 988 3123 992
rect 279 968 343 972
rect 2969 968 3033 972
rect 369 878 433 882
rect 3059 878 3123 882
rect 279 858 343 862
rect 2969 858 3033 862
rect 369 768 433 772
rect 1624 767 1628 771
rect 3059 768 3123 772
rect 1664 757 1668 761
rect 1672 757 1676 761
rect 279 748 343 752
rect 2969 748 3033 752
rect 1656 693 1660 697
rect 1664 693 1668 697
rect 369 658 433 662
rect 1624 657 1628 661
rect 3059 658 3123 662
rect 1664 647 1668 651
rect 1672 647 1676 651
rect 279 638 343 642
rect 2969 638 3033 642
rect 712 592 716 596
rect 1656 583 1660 587
rect 1664 583 1668 587
rect 369 548 433 552
rect 1624 547 1628 551
rect 3059 548 3123 552
rect 1664 537 1668 541
rect 1672 537 1676 541
rect 279 528 343 532
rect 2969 528 3033 532
rect 720 482 724 486
rect 1656 473 1660 477
rect 1664 473 1668 477
rect 369 438 433 442
rect 1624 437 1628 441
rect 3059 438 3123 442
rect 1664 427 1668 431
rect 1672 427 1676 431
rect 279 418 343 422
rect 2969 418 3033 422
rect 728 372 732 376
rect 1656 363 1660 367
rect 1664 363 1668 367
rect 2216 363 2220 367
rect 369 328 433 332
rect 1624 327 1628 331
rect 3059 328 3123 332
rect 1664 317 1668 321
rect 1672 317 1676 321
rect 279 308 343 312
rect 2969 308 3033 312
rect 736 262 740 266
rect 1656 253 1660 257
rect 1664 253 1668 257
rect 369 218 433 222
rect 1624 217 1628 221
rect 3059 218 3123 222
rect 1664 207 1668 211
rect 1672 207 1676 211
rect 279 198 343 202
rect 2969 198 3033 202
rect 744 152 748 156
rect 369 108 433 112
rect 1624 107 1628 111
rect 1672 107 1676 111
rect 3059 108 3123 112
rect 279 88 343 92
rect 1624 87 1628 91
rect 2969 88 3033 92
rect 752 42 756 46
rect 1656 33 1660 37
rect 1664 33 1668 37
rect 369 -2 433 2
rect 1672 -3 1676 1
rect 3059 -2 3123 2
<< metal2 >>
rect 279 1302 343 1343
rect 279 1192 343 1298
rect 279 1082 343 1188
rect 279 972 343 1078
rect 279 862 343 968
rect 279 752 343 858
rect 279 642 343 748
rect 279 532 343 638
rect 279 422 343 528
rect 279 312 343 418
rect 279 202 343 308
rect 279 92 343 198
rect 279 58 343 88
rect 369 1212 433 1342
rect 369 1102 433 1208
rect 369 992 433 1098
rect 369 882 433 988
rect 369 772 433 878
rect 369 662 433 768
rect 369 552 433 658
rect 369 442 433 548
rect 369 332 433 438
rect 369 222 433 328
rect 369 112 433 218
rect 369 2 433 108
rect 462 82 466 1577
rect 469 192 473 1687
rect 476 302 480 1797
rect 483 412 487 1907
rect 490 522 494 2017
rect 497 632 501 2127
rect 504 742 508 2237
rect 512 852 516 2347
rect 520 918 524 1312
rect 544 1202 548 1312
rect 552 1222 556 1312
rect 559 962 563 2457
rect 566 952 570 2447
rect 582 2417 586 2811
rect 661 2741 667 2742
rect 661 2737 662 2741
rect 666 2737 667 2741
rect 661 2736 667 2737
rect 662 2462 666 2736
rect 661 2461 667 2462
rect 661 2457 662 2461
rect 666 2457 667 2461
rect 661 2456 667 2457
rect 613 2451 619 2452
rect 613 2447 614 2451
rect 618 2447 619 2451
rect 613 2446 619 2447
rect 614 2438 618 2446
rect 662 2438 666 2456
rect 589 2351 595 2352
rect 589 2347 590 2351
rect 594 2347 595 2351
rect 589 2346 595 2347
rect 590 2312 594 2346
rect 710 2315 714 2811
rect 589 2241 595 2242
rect 589 2237 590 2241
rect 594 2237 595 2241
rect 589 2236 595 2237
rect 590 2202 594 2236
rect 718 2205 722 2811
rect 589 2131 595 2132
rect 589 2127 590 2131
rect 594 2127 595 2131
rect 589 2126 595 2127
rect 590 2092 594 2126
rect 726 2095 730 2811
rect 589 2021 595 2022
rect 589 2017 590 2021
rect 594 2017 595 2021
rect 589 2016 595 2017
rect 590 1982 594 2016
rect 734 1985 738 2811
rect 589 1911 595 1912
rect 589 1907 590 1911
rect 594 1907 595 1911
rect 589 1906 595 1907
rect 590 1872 594 1906
rect 742 1875 746 2811
rect 589 1801 595 1802
rect 589 1797 590 1801
rect 594 1797 595 1801
rect 589 1796 595 1797
rect 590 1762 594 1796
rect 750 1765 754 2811
rect 766 2417 770 2811
rect 845 2461 851 2462
rect 845 2457 846 2461
rect 850 2457 851 2461
rect 845 2456 851 2457
rect 797 2451 803 2452
rect 797 2447 798 2451
rect 802 2447 803 2451
rect 797 2446 803 2447
rect 798 2438 802 2446
rect 846 2438 850 2456
rect 950 2417 954 2811
rect 1029 2461 1035 2462
rect 1029 2457 1030 2461
rect 1034 2457 1035 2461
rect 1029 2456 1035 2457
rect 981 2451 987 2452
rect 981 2447 982 2451
rect 986 2447 987 2451
rect 981 2446 987 2447
rect 982 2438 986 2446
rect 1030 2438 1034 2456
rect 773 2351 779 2352
rect 773 2347 774 2351
rect 778 2347 779 2351
rect 773 2346 779 2347
rect 957 2351 963 2352
rect 957 2347 958 2351
rect 962 2347 963 2351
rect 957 2346 963 2347
rect 774 2312 778 2346
rect 958 2312 962 2346
rect 773 2241 779 2242
rect 773 2237 774 2241
rect 778 2237 779 2241
rect 773 2236 779 2237
rect 774 2202 778 2236
rect 773 2131 779 2132
rect 773 2127 774 2131
rect 778 2127 779 2131
rect 773 2126 779 2127
rect 774 2092 778 2126
rect 773 2021 779 2022
rect 773 2017 774 2021
rect 778 2017 779 2021
rect 773 2016 779 2017
rect 774 1982 778 2016
rect 773 1911 779 1912
rect 773 1907 774 1911
rect 778 1907 779 1911
rect 773 1906 779 1907
rect 774 1872 778 1906
rect 773 1801 779 1802
rect 773 1797 774 1801
rect 778 1797 779 1801
rect 773 1796 779 1797
rect 774 1762 778 1796
rect 589 1691 595 1692
rect 589 1687 590 1691
rect 594 1687 595 1691
rect 589 1686 595 1687
rect 773 1691 779 1692
rect 773 1687 774 1691
rect 778 1687 779 1691
rect 773 1686 779 1687
rect 590 1652 594 1686
rect 774 1652 778 1686
rect 589 1581 595 1582
rect 589 1577 590 1581
rect 594 1577 595 1581
rect 589 1576 595 1577
rect 773 1581 779 1582
rect 773 1577 774 1581
rect 778 1577 779 1581
rect 773 1576 779 1577
rect 590 1542 594 1576
rect 774 1542 778 1576
rect 584 918 588 1312
rect 615 1222 621 1223
rect 615 1218 616 1222
rect 620 1218 621 1222
rect 615 1217 621 1218
rect 616 953 620 1217
rect 636 1042 640 1481
rect 643 1152 647 1471
rect 650 1262 654 1460
rect 657 1182 661 1450
rect 657 1062 661 1178
rect 665 1172 669 1440
rect 665 1162 669 1168
rect 672 1282 676 1430
rect 672 1132 676 1278
rect 680 1072 684 1420
rect 688 1052 692 1410
rect 894 1403 898 2311
rect 957 2241 963 2242
rect 957 2237 958 2241
rect 962 2237 963 2241
rect 957 2236 963 2237
rect 958 2202 962 2236
rect 902 1414 906 2201
rect 957 2131 963 2132
rect 957 2127 958 2131
rect 962 2127 963 2131
rect 957 2126 963 2127
rect 958 2092 962 2126
rect 910 1424 914 2091
rect 957 2021 963 2022
rect 957 2017 958 2021
rect 962 2017 963 2021
rect 957 2016 963 2017
rect 958 1982 962 2016
rect 957 1911 963 1912
rect 957 1907 958 1911
rect 962 1907 963 1911
rect 957 1906 963 1907
rect 958 1872 962 1906
rect 957 1801 963 1802
rect 957 1797 958 1801
rect 962 1797 963 1801
rect 957 1796 963 1797
rect 958 1762 962 1796
rect 918 1434 922 1761
rect 957 1691 963 1692
rect 957 1687 958 1691
rect 962 1687 963 1691
rect 957 1686 963 1687
rect 958 1652 962 1686
rect 926 1444 930 1651
rect 957 1581 963 1582
rect 957 1577 958 1581
rect 962 1577 963 1581
rect 957 1576 963 1577
rect 958 1542 962 1576
rect 934 1454 938 1541
rect 1078 1464 1082 2091
rect 1086 1475 1090 1981
rect 1094 1485 1098 1871
rect 663 962 669 963
rect 663 958 664 962
rect 668 958 669 962
rect 663 957 669 958
rect 615 952 621 953
rect 615 948 616 952
rect 620 948 621 952
rect 615 947 621 948
rect 616 939 620 947
rect 664 939 668 957
rect 696 943 700 1388
rect 704 1022 708 1399
rect 695 942 701 943
rect 695 938 696 942
rect 700 938 701 942
rect 695 937 701 938
rect 591 852 597 853
rect 591 848 592 852
rect 596 848 597 852
rect 591 847 597 848
rect 559 832 565 833
rect 559 828 560 832
rect 564 828 565 832
rect 559 827 565 828
rect 520 813 524 819
rect 519 812 525 813
rect 519 808 520 812
rect 524 808 525 812
rect 519 807 525 808
rect 552 803 556 818
rect 560 808 564 827
rect 592 813 596 847
rect 703 832 709 833
rect 703 828 704 832
rect 708 828 709 832
rect 703 827 709 828
rect 704 812 708 827
rect 551 802 557 803
rect 551 798 552 802
rect 556 798 557 802
rect 551 797 557 798
rect 591 742 597 743
rect 591 738 592 742
rect 596 738 597 742
rect 591 737 597 738
rect 559 722 565 723
rect 559 718 560 722
rect 564 718 565 722
rect 559 717 565 718
rect 520 703 524 709
rect 519 702 525 703
rect 519 698 520 702
rect 524 698 525 702
rect 519 697 525 698
rect 552 693 556 708
rect 560 698 564 717
rect 592 703 596 737
rect 703 722 709 723
rect 703 718 704 722
rect 708 718 709 722
rect 703 717 709 718
rect 704 702 708 717
rect 551 692 557 693
rect 551 688 552 692
rect 556 688 557 692
rect 551 687 557 688
rect 591 632 597 633
rect 591 628 592 632
rect 596 628 597 632
rect 591 627 597 628
rect 559 612 565 613
rect 559 608 560 612
rect 564 608 565 612
rect 559 607 565 608
rect 520 593 524 599
rect 519 592 525 593
rect 519 588 520 592
rect 524 588 525 592
rect 519 587 525 588
rect 552 583 556 598
rect 560 588 564 607
rect 592 593 596 627
rect 703 612 709 613
rect 703 608 704 612
rect 708 608 709 612
rect 703 607 709 608
rect 704 592 708 607
rect 712 596 716 1378
rect 551 582 557 583
rect 551 578 552 582
rect 556 578 557 582
rect 551 577 557 578
rect 591 522 597 523
rect 591 518 592 522
rect 596 518 597 522
rect 591 517 597 518
rect 559 502 565 503
rect 559 498 560 502
rect 564 498 565 502
rect 559 497 565 498
rect 520 483 524 489
rect 519 482 525 483
rect 519 478 520 482
rect 524 478 525 482
rect 519 477 525 478
rect 552 473 556 488
rect 560 478 564 497
rect 592 483 596 517
rect 703 502 709 503
rect 703 498 704 502
rect 708 498 709 502
rect 703 497 709 498
rect 704 482 708 497
rect 720 486 724 1368
rect 551 472 557 473
rect 551 468 552 472
rect 556 468 557 472
rect 551 467 557 468
rect 591 412 597 413
rect 591 408 592 412
rect 596 408 597 412
rect 591 407 597 408
rect 559 392 565 393
rect 559 388 560 392
rect 564 388 565 392
rect 559 387 565 388
rect 520 373 524 379
rect 519 372 525 373
rect 519 368 520 372
rect 524 368 525 372
rect 519 367 525 368
rect 552 363 556 378
rect 560 368 564 387
rect 592 373 596 407
rect 703 392 709 393
rect 703 388 704 392
rect 708 388 709 392
rect 703 387 709 388
rect 704 372 708 387
rect 728 376 732 1358
rect 551 362 557 363
rect 551 358 552 362
rect 556 358 557 362
rect 551 357 557 358
rect 591 302 597 303
rect 591 298 592 302
rect 596 298 597 302
rect 591 297 597 298
rect 559 282 565 283
rect 559 278 560 282
rect 564 278 565 282
rect 559 277 565 278
rect 520 263 524 269
rect 519 262 525 263
rect 519 258 520 262
rect 524 258 525 262
rect 519 257 525 258
rect 552 253 556 268
rect 560 258 564 277
rect 592 263 596 297
rect 703 282 709 283
rect 703 278 704 282
rect 708 278 709 282
rect 703 277 709 278
rect 704 262 708 277
rect 736 266 740 1348
rect 551 252 557 253
rect 551 248 552 252
rect 556 248 557 252
rect 551 247 557 248
rect 591 192 597 193
rect 591 188 592 192
rect 596 188 597 192
rect 591 187 597 188
rect 559 172 565 173
rect 559 168 560 172
rect 564 168 565 172
rect 559 167 565 168
rect 520 153 524 159
rect 519 152 525 153
rect 519 148 520 152
rect 524 148 525 152
rect 519 147 525 148
rect 552 143 556 158
rect 560 148 564 167
rect 592 153 596 187
rect 703 172 709 173
rect 703 168 704 172
rect 708 168 709 172
rect 703 167 709 168
rect 704 152 708 167
rect 744 156 748 1338
rect 551 142 557 143
rect 551 138 552 142
rect 556 138 557 142
rect 551 137 557 138
rect 591 82 597 83
rect 591 78 592 82
rect 596 78 597 82
rect 591 77 597 78
rect 559 62 565 63
rect 559 58 560 62
rect 564 58 565 62
rect 559 57 565 58
rect 520 43 524 49
rect 519 42 525 43
rect 519 38 520 42
rect 524 38 525 42
rect 519 37 525 38
rect 552 33 556 48
rect 560 38 564 57
rect 592 43 596 77
rect 703 62 709 63
rect 703 58 704 62
rect 708 58 709 62
rect 703 57 709 58
rect 704 42 708 57
rect 752 46 756 1328
rect 767 1262 773 1263
rect 767 1258 768 1262
rect 772 1258 773 1262
rect 767 1257 773 1258
rect 768 1254 772 1257
rect 767 1152 773 1153
rect 767 1148 768 1152
rect 772 1148 773 1152
rect 767 1147 773 1148
rect 768 1144 772 1147
rect 767 1042 773 1043
rect 767 1038 768 1042
rect 772 1038 773 1042
rect 792 1041 796 1318
rect 799 1282 805 1283
rect 799 1278 800 1282
rect 804 1278 805 1282
rect 799 1277 805 1278
rect 800 1264 804 1277
rect 856 1202 860 1251
rect 888 1202 892 1251
rect 960 1248 964 1308
rect 799 1172 805 1173
rect 799 1168 800 1172
rect 804 1168 805 1172
rect 799 1167 805 1168
rect 800 1154 804 1167
rect 816 1139 820 1198
rect 872 1092 876 1198
rect 799 1062 805 1063
rect 799 1058 800 1062
rect 804 1058 805 1062
rect 799 1057 805 1058
rect 800 1044 804 1057
rect 767 1037 773 1038
rect 768 1034 772 1037
rect 816 1029 820 1088
rect 815 962 821 963
rect 815 958 816 962
rect 820 958 821 962
rect 815 957 821 958
rect 1551 962 1557 963
rect 1551 958 1552 962
rect 1556 958 1557 962
rect 1551 957 1557 958
rect 767 952 773 953
rect 767 948 768 952
rect 772 948 773 952
rect 767 947 773 948
rect 768 939 772 947
rect 816 939 820 957
rect 1503 952 1509 953
rect 1503 948 1504 952
rect 1508 948 1509 952
rect 1503 947 1509 948
rect 871 942 877 943
rect 871 938 872 942
rect 876 938 877 942
rect 1504 939 1508 947
rect 1552 939 1556 957
rect 871 937 877 938
rect 872 919 876 937
rect 1600 918 1604 1312
rect 1632 918 1636 1312
rect 1670 872 1674 1036
rect 767 852 773 853
rect 767 848 768 852
rect 772 848 773 852
rect 767 847 773 848
rect 768 813 772 847
rect 1591 842 1597 843
rect 1591 838 1592 842
rect 1596 838 1597 842
rect 1591 837 1597 838
rect 1615 842 1621 843
rect 1615 838 1616 842
rect 1620 838 1621 842
rect 1615 837 1621 838
rect 911 822 917 823
rect 911 818 912 822
rect 916 818 917 822
rect 911 817 917 818
rect 904 813 908 817
rect 903 812 909 813
rect 903 808 904 812
rect 908 808 909 812
rect 912 809 916 817
rect 903 807 909 808
rect 1504 783 1508 816
rect 1592 812 1596 837
rect 1616 804 1620 837
rect 1656 833 1660 868
rect 1655 832 1661 833
rect 1655 828 1656 832
rect 1660 828 1661 832
rect 1655 827 1661 828
rect 1671 832 1677 833
rect 1671 828 1672 832
rect 1676 828 1677 832
rect 1671 827 1677 828
rect 1656 819 1660 827
rect 1503 782 1509 783
rect 1503 778 1504 782
rect 1508 778 1509 782
rect 1503 777 1509 778
rect 1624 771 1628 807
rect 1672 761 1676 827
rect 767 742 773 743
rect 767 738 768 742
rect 772 738 773 742
rect 767 737 773 738
rect 768 703 772 737
rect 1591 732 1597 733
rect 1591 728 1592 732
rect 1596 728 1597 732
rect 1591 727 1597 728
rect 1615 732 1621 733
rect 1615 728 1616 732
rect 1620 728 1621 732
rect 1615 727 1621 728
rect 911 712 917 713
rect 911 708 912 712
rect 916 708 917 712
rect 911 707 917 708
rect 904 703 908 707
rect 903 702 909 703
rect 903 698 904 702
rect 908 698 909 702
rect 912 699 916 707
rect 903 697 909 698
rect 1504 673 1508 706
rect 1592 702 1596 727
rect 1616 694 1620 727
rect 1624 722 1628 759
rect 1688 763 1692 1036
rect 1759 962 1765 963
rect 1759 958 1760 962
rect 1764 958 1765 962
rect 1759 957 1765 958
rect 1711 952 1717 953
rect 1711 948 1712 952
rect 1716 948 1717 952
rect 1711 947 1717 948
rect 1712 939 1716 947
rect 1760 939 1764 957
rect 1808 918 1812 1312
rect 1911 962 1917 963
rect 1911 958 1912 962
rect 1916 958 1917 962
rect 1911 957 1917 958
rect 1863 952 1869 953
rect 1863 948 1864 952
rect 1868 948 1869 952
rect 1863 947 1869 948
rect 1864 939 1868 947
rect 1912 939 1916 957
rect 1960 918 1964 1312
rect 1992 918 1996 1312
rect 2048 918 2052 1312
rect 2079 1202 2085 1203
rect 2079 1198 2080 1202
rect 2084 1198 2085 1202
rect 2079 1197 2085 1198
rect 2080 918 2084 1197
rect 2143 962 2149 963
rect 2143 958 2144 962
rect 2148 958 2149 962
rect 2143 957 2149 958
rect 2095 952 2101 953
rect 2095 948 2096 952
rect 2100 948 2101 952
rect 2095 947 2101 948
rect 2096 939 2100 947
rect 2144 939 2148 957
rect 1847 851 1853 852
rect 1847 847 1848 851
rect 1852 847 1853 851
rect 1847 846 1853 847
rect 1695 842 1701 843
rect 1695 838 1696 842
rect 1700 838 1701 842
rect 1695 837 1701 838
rect 1696 807 1700 837
rect 1712 793 1716 816
rect 1840 803 1844 818
rect 1848 808 1852 846
rect 2015 832 2021 833
rect 2015 828 2016 832
rect 2020 828 2021 832
rect 2015 827 2021 828
rect 1839 802 1845 803
rect 1839 798 1840 802
rect 1844 798 1845 802
rect 1839 797 1845 798
rect 1711 792 1717 793
rect 1711 788 1712 792
rect 1716 788 1717 792
rect 1711 787 1717 788
rect 1864 783 1868 816
rect 1952 813 1956 815
rect 1976 813 1980 821
rect 2016 818 2020 827
rect 1951 812 1957 813
rect 1975 812 1981 813
rect 1951 808 1952 812
rect 1956 808 1957 812
rect 1951 807 1957 808
rect 1968 783 1972 812
rect 1975 808 1976 812
rect 1980 808 1981 812
rect 1975 807 1981 808
rect 2176 803 2180 812
rect 2175 802 2181 803
rect 2175 798 2176 802
rect 2180 798 2181 802
rect 2175 797 2181 798
rect 1863 782 1869 783
rect 1863 778 1864 782
rect 1868 778 1869 782
rect 1863 777 1869 778
rect 1967 782 1973 783
rect 1967 778 1968 782
rect 1972 778 1973 782
rect 1967 777 1973 778
rect 1655 722 1661 723
rect 1655 718 1656 722
rect 1660 718 1661 722
rect 1655 717 1661 718
rect 1656 709 1660 717
rect 1664 697 1668 757
rect 1847 741 1853 742
rect 1847 737 1848 741
rect 1852 737 1853 741
rect 1847 736 1853 737
rect 1695 732 1701 733
rect 1695 728 1696 732
rect 1700 728 1701 732
rect 1695 727 1701 728
rect 1671 722 1677 723
rect 1671 718 1672 722
rect 1676 718 1677 722
rect 1671 717 1677 718
rect 1503 672 1509 673
rect 1503 668 1504 672
rect 1508 668 1509 672
rect 1503 667 1509 668
rect 1624 661 1628 697
rect 767 632 773 633
rect 767 628 768 632
rect 772 628 773 632
rect 767 627 773 628
rect 768 593 772 627
rect 1591 622 1597 623
rect 1591 618 1592 622
rect 1596 618 1597 622
rect 1591 617 1597 618
rect 1615 622 1621 623
rect 1615 618 1616 622
rect 1620 618 1621 622
rect 1615 617 1621 618
rect 911 602 917 603
rect 911 598 912 602
rect 916 598 917 602
rect 911 597 917 598
rect 904 593 908 597
rect 903 592 909 593
rect 903 588 904 592
rect 908 588 909 592
rect 912 589 916 597
rect 903 587 909 588
rect 1504 563 1508 596
rect 1592 592 1596 617
rect 1616 584 1620 617
rect 1656 613 1660 693
rect 1672 651 1676 717
rect 1696 697 1700 727
rect 1712 683 1716 706
rect 1840 693 1844 708
rect 1848 698 1852 736
rect 2015 722 2021 723
rect 2015 718 2016 722
rect 2020 718 2021 722
rect 2015 717 2021 718
rect 1839 692 1845 693
rect 1839 688 1840 692
rect 1844 688 1845 692
rect 1839 687 1845 688
rect 1711 682 1717 683
rect 1711 678 1712 682
rect 1716 678 1717 682
rect 1711 677 1717 678
rect 1864 673 1868 706
rect 1952 703 1956 705
rect 1976 703 1980 711
rect 2016 708 2020 717
rect 1951 702 1957 703
rect 1975 702 1981 703
rect 1951 698 1952 702
rect 1956 698 1957 702
rect 1951 697 1957 698
rect 1968 673 1972 702
rect 1975 698 1976 702
rect 1980 698 1981 702
rect 1975 697 1981 698
rect 2176 693 2180 702
rect 2175 692 2181 693
rect 2175 688 2176 692
rect 2180 688 2181 692
rect 2175 687 2181 688
rect 1863 672 1869 673
rect 1863 668 1864 672
rect 1868 668 1869 672
rect 1863 667 1869 668
rect 1967 672 1973 673
rect 1967 668 1968 672
rect 1972 668 1973 672
rect 1967 667 1973 668
rect 1655 612 1661 613
rect 1655 608 1656 612
rect 1660 608 1661 612
rect 1655 607 1661 608
rect 1656 599 1660 607
rect 1664 587 1668 647
rect 1847 631 1853 632
rect 1847 627 1848 631
rect 1852 627 1853 631
rect 1847 626 1853 627
rect 1695 622 1701 623
rect 1695 618 1696 622
rect 1700 618 1701 622
rect 1695 617 1701 618
rect 1671 612 1677 613
rect 1671 608 1672 612
rect 1676 608 1677 612
rect 1671 607 1677 608
rect 1503 562 1509 563
rect 1503 558 1504 562
rect 1508 558 1509 562
rect 1503 557 1509 558
rect 1624 551 1628 587
rect 767 522 773 523
rect 767 518 768 522
rect 772 518 773 522
rect 767 517 773 518
rect 768 483 772 517
rect 1591 512 1597 513
rect 1591 508 1592 512
rect 1596 508 1597 512
rect 1591 507 1597 508
rect 1615 512 1621 513
rect 1615 508 1616 512
rect 1620 508 1621 512
rect 1615 507 1621 508
rect 911 492 917 493
rect 911 488 912 492
rect 916 488 917 492
rect 911 487 917 488
rect 904 483 908 487
rect 903 482 909 483
rect 903 478 904 482
rect 908 478 909 482
rect 912 479 916 487
rect 903 477 909 478
rect 1504 453 1508 486
rect 1592 482 1596 507
rect 1616 474 1620 507
rect 1656 503 1660 583
rect 1672 541 1676 607
rect 1696 587 1700 617
rect 1712 573 1716 596
rect 1840 583 1844 598
rect 1848 588 1852 626
rect 2015 612 2021 613
rect 2015 608 2016 612
rect 2020 608 2021 612
rect 2015 607 2021 608
rect 1839 582 1845 583
rect 1839 578 1840 582
rect 1844 578 1845 582
rect 1839 577 1845 578
rect 1711 572 1717 573
rect 1711 568 1712 572
rect 1716 568 1717 572
rect 1711 567 1717 568
rect 1864 563 1868 596
rect 1952 593 1956 595
rect 1976 593 1980 601
rect 2016 598 2020 607
rect 1951 592 1957 593
rect 1975 592 1981 593
rect 1951 588 1952 592
rect 1956 588 1957 592
rect 1951 587 1957 588
rect 1968 563 1972 592
rect 1975 588 1976 592
rect 1980 588 1981 592
rect 1975 587 1981 588
rect 2176 583 2180 592
rect 2175 582 2181 583
rect 2175 578 2176 582
rect 2180 578 2181 582
rect 2175 577 2181 578
rect 1863 562 1869 563
rect 1863 558 1864 562
rect 1868 558 1869 562
rect 1863 557 1869 558
rect 1967 562 1973 563
rect 1967 558 1968 562
rect 1972 558 1973 562
rect 1967 557 1973 558
rect 1655 502 1661 503
rect 1655 498 1656 502
rect 1660 498 1661 502
rect 1655 497 1661 498
rect 1656 489 1660 497
rect 1664 477 1668 537
rect 1847 521 1853 522
rect 1847 517 1848 521
rect 1852 517 1853 521
rect 1847 516 1853 517
rect 1695 512 1701 513
rect 1695 508 1696 512
rect 1700 508 1701 512
rect 1695 507 1701 508
rect 1671 502 1677 503
rect 1671 498 1672 502
rect 1676 498 1677 502
rect 1671 497 1677 498
rect 1503 452 1509 453
rect 1503 448 1504 452
rect 1508 448 1509 452
rect 1503 447 1509 448
rect 1624 441 1628 477
rect 767 412 773 413
rect 767 408 768 412
rect 772 408 773 412
rect 767 407 773 408
rect 768 373 772 407
rect 1591 402 1597 403
rect 1591 398 1592 402
rect 1596 398 1597 402
rect 1591 397 1597 398
rect 1615 402 1621 403
rect 1615 398 1616 402
rect 1620 398 1621 402
rect 1615 397 1621 398
rect 911 382 917 383
rect 911 378 912 382
rect 916 378 917 382
rect 911 377 917 378
rect 904 373 908 377
rect 903 372 909 373
rect 903 368 904 372
rect 908 368 909 372
rect 912 369 916 377
rect 903 367 909 368
rect 1504 343 1508 376
rect 1592 372 1596 397
rect 1616 364 1620 397
rect 1656 393 1660 473
rect 1672 431 1676 497
rect 1696 477 1700 507
rect 1712 463 1716 486
rect 1840 473 1844 488
rect 1848 478 1852 516
rect 2015 502 2021 503
rect 2015 498 2016 502
rect 2020 498 2021 502
rect 2015 497 2021 498
rect 1839 472 1845 473
rect 1839 468 1840 472
rect 1844 468 1845 472
rect 1839 467 1845 468
rect 1711 462 1717 463
rect 1711 458 1712 462
rect 1716 458 1717 462
rect 1711 457 1717 458
rect 1864 453 1868 486
rect 1952 483 1956 485
rect 1976 483 1980 491
rect 2016 488 2020 497
rect 1951 482 1957 483
rect 1975 482 1981 483
rect 1951 478 1952 482
rect 1956 478 1957 482
rect 1951 477 1957 478
rect 1968 453 1972 482
rect 1975 478 1976 482
rect 1980 478 1981 482
rect 1975 477 1981 478
rect 2176 473 2180 482
rect 2175 472 2181 473
rect 2175 468 2176 472
rect 2180 468 2181 472
rect 2175 467 2181 468
rect 1863 452 1869 453
rect 1863 448 1864 452
rect 1868 448 1869 452
rect 1863 447 1869 448
rect 1967 452 1973 453
rect 1967 448 1968 452
rect 1972 448 1973 452
rect 1967 447 1973 448
rect 1655 392 1661 393
rect 1655 388 1656 392
rect 1660 388 1661 392
rect 1655 387 1661 388
rect 1656 379 1660 387
rect 1664 367 1668 427
rect 1847 411 1853 412
rect 1847 407 1848 411
rect 1852 407 1853 411
rect 1847 406 1853 407
rect 1695 402 1701 403
rect 1695 398 1696 402
rect 1700 398 1701 402
rect 1695 397 1701 398
rect 1671 392 1677 393
rect 1671 388 1672 392
rect 1676 388 1677 392
rect 1671 387 1677 388
rect 1503 342 1509 343
rect 1503 338 1504 342
rect 1508 338 1509 342
rect 1503 337 1509 338
rect 1624 331 1628 367
rect 767 302 773 303
rect 767 298 768 302
rect 772 298 773 302
rect 767 297 773 298
rect 768 263 772 297
rect 1591 292 1597 293
rect 1591 288 1592 292
rect 1596 288 1597 292
rect 1591 287 1597 288
rect 1615 292 1621 293
rect 1615 288 1616 292
rect 1620 288 1621 292
rect 1615 287 1621 288
rect 911 272 917 273
rect 911 268 912 272
rect 916 268 917 272
rect 911 267 917 268
rect 904 263 908 267
rect 903 262 909 263
rect 903 258 904 262
rect 908 258 909 262
rect 912 259 916 267
rect 903 257 909 258
rect 1504 233 1508 266
rect 1592 262 1596 287
rect 1616 254 1620 287
rect 1656 283 1660 363
rect 1672 321 1676 387
rect 1696 367 1700 397
rect 1712 353 1716 376
rect 1840 363 1844 378
rect 1848 368 1852 406
rect 2015 392 2021 393
rect 2015 388 2016 392
rect 2020 388 2021 392
rect 2015 387 2021 388
rect 1839 362 1845 363
rect 1839 358 1840 362
rect 1844 358 1845 362
rect 1839 357 1845 358
rect 1711 352 1717 353
rect 1711 348 1712 352
rect 1716 348 1717 352
rect 1711 347 1717 348
rect 1864 343 1868 376
rect 1952 373 1956 375
rect 1976 373 1980 381
rect 2016 378 2020 387
rect 1951 372 1957 373
rect 1975 372 1981 373
rect 1951 368 1952 372
rect 1956 368 1957 372
rect 1951 367 1957 368
rect 1968 343 1972 372
rect 1975 368 1976 372
rect 1980 368 1981 372
rect 1975 367 1981 368
rect 2176 363 2180 372
rect 2216 367 2220 1312
rect 2271 884 2275 1312
rect 2279 884 2283 1312
rect 2311 884 2315 1312
rect 2327 884 2331 1312
rect 2344 884 2348 1312
rect 2463 982 2467 1312
rect 2503 982 2507 1312
rect 2807 1310 2811 1314
rect 2969 1302 3033 1343
rect 2969 1192 3033 1298
rect 2871 1092 2875 1096
rect 2969 1082 3033 1188
rect 2919 984 2923 988
rect 2969 972 3033 1078
rect 2969 862 3033 968
rect 2969 752 3033 858
rect 2969 642 3033 748
rect 2969 532 3033 638
rect 2969 422 3033 528
rect 2175 362 2181 363
rect 2175 358 2176 362
rect 2180 358 2181 362
rect 2175 357 2181 358
rect 1863 342 1869 343
rect 1863 338 1864 342
rect 1868 338 1869 342
rect 1863 337 1869 338
rect 1967 342 1973 343
rect 1967 338 1968 342
rect 1972 338 1973 342
rect 1967 337 1973 338
rect 1655 282 1661 283
rect 1655 278 1656 282
rect 1660 278 1661 282
rect 1655 277 1661 278
rect 1656 269 1660 277
rect 1664 257 1668 317
rect 2969 312 3033 418
rect 1847 301 1853 302
rect 1847 297 1848 301
rect 1852 297 1853 301
rect 1847 296 1853 297
rect 1695 292 1701 293
rect 1695 288 1696 292
rect 1700 288 1701 292
rect 1695 287 1701 288
rect 1671 282 1677 283
rect 1671 278 1672 282
rect 1676 278 1677 282
rect 1671 277 1677 278
rect 1503 232 1509 233
rect 1503 228 1504 232
rect 1508 228 1509 232
rect 1503 227 1509 228
rect 1624 221 1628 257
rect 767 192 773 193
rect 767 188 768 192
rect 772 188 773 192
rect 767 187 773 188
rect 768 153 772 187
rect 1591 182 1597 183
rect 1591 178 1592 182
rect 1596 178 1597 182
rect 1591 177 1597 178
rect 1615 182 1621 183
rect 1615 178 1616 182
rect 1620 178 1621 182
rect 1615 177 1621 178
rect 911 162 917 163
rect 911 158 912 162
rect 916 158 917 162
rect 911 157 917 158
rect 904 153 908 157
rect 903 152 909 153
rect 903 148 904 152
rect 908 148 909 152
rect 912 149 916 157
rect 903 147 909 148
rect 1504 123 1508 156
rect 1592 152 1596 177
rect 1616 144 1620 177
rect 1656 173 1660 253
rect 1672 211 1676 277
rect 1696 257 1700 287
rect 1712 243 1716 266
rect 1840 253 1844 268
rect 1848 258 1852 296
rect 2015 282 2021 283
rect 2015 278 2016 282
rect 2020 278 2021 282
rect 2015 277 2021 278
rect 1839 252 1845 253
rect 1839 248 1840 252
rect 1844 248 1845 252
rect 1839 247 1845 248
rect 1711 242 1717 243
rect 1711 238 1712 242
rect 1716 238 1717 242
rect 1711 237 1717 238
rect 1864 233 1868 266
rect 1952 263 1956 265
rect 1976 263 1980 271
rect 2016 268 2020 277
rect 1951 262 1957 263
rect 1975 262 1981 263
rect 1951 258 1952 262
rect 1956 258 1957 262
rect 1951 257 1957 258
rect 1968 233 1972 262
rect 1975 258 1976 262
rect 1980 258 1981 262
rect 1975 257 1981 258
rect 2176 253 2180 262
rect 2175 252 2181 253
rect 2175 248 2176 252
rect 2180 248 2181 252
rect 2175 247 2181 248
rect 1863 232 1869 233
rect 1863 228 1864 232
rect 1868 228 1869 232
rect 1863 227 1869 228
rect 1967 232 1973 233
rect 1967 228 1968 232
rect 1972 228 1973 232
rect 1967 227 1973 228
rect 1655 172 1661 173
rect 1655 168 1656 172
rect 1660 168 1661 172
rect 1655 167 1661 168
rect 1656 159 1660 167
rect 1503 122 1509 123
rect 1503 118 1504 122
rect 1508 118 1509 122
rect 1503 117 1509 118
rect 1624 111 1628 147
rect 767 82 773 83
rect 767 78 768 82
rect 772 78 773 82
rect 767 77 773 78
rect 768 43 772 77
rect 1591 72 1597 73
rect 1591 68 1592 72
rect 1596 68 1597 72
rect 1591 67 1597 68
rect 1615 72 1621 73
rect 1615 68 1616 72
rect 1620 68 1621 72
rect 1615 67 1621 68
rect 911 52 917 53
rect 911 48 912 52
rect 916 48 917 52
rect 911 47 917 48
rect 904 43 908 47
rect 903 42 909 43
rect 903 38 904 42
rect 908 38 909 42
rect 912 39 916 47
rect 903 37 909 38
rect 551 32 557 33
rect 551 28 552 32
rect 556 28 557 32
rect 551 27 557 28
rect 1504 13 1508 46
rect 1592 42 1596 67
rect 1616 34 1620 67
rect 1624 34 1628 87
rect 1655 62 1661 63
rect 1655 58 1656 62
rect 1660 58 1661 62
rect 1655 57 1661 58
rect 1656 37 1660 57
rect 1664 37 1668 207
rect 2969 202 3033 308
rect 1847 191 1853 192
rect 1847 187 1848 191
rect 1852 187 1853 191
rect 1847 186 1853 187
rect 1695 182 1701 183
rect 1695 178 1696 182
rect 1700 178 1701 182
rect 1695 177 1701 178
rect 1671 172 1677 173
rect 1671 168 1672 172
rect 1676 168 1677 172
rect 1671 167 1677 168
rect 1672 111 1676 167
rect 1696 147 1700 177
rect 1712 133 1716 156
rect 1840 143 1844 158
rect 1848 148 1852 186
rect 2015 172 2021 173
rect 2015 168 2016 172
rect 2020 168 2021 172
rect 2015 167 2021 168
rect 1839 142 1845 143
rect 1839 138 1840 142
rect 1844 138 1845 142
rect 1839 137 1845 138
rect 1711 132 1717 133
rect 1711 128 1712 132
rect 1716 128 1717 132
rect 1711 127 1717 128
rect 1864 123 1868 156
rect 1952 153 1956 155
rect 1976 153 1980 161
rect 2016 158 2020 167
rect 1951 152 1957 153
rect 1975 152 1981 153
rect 1951 148 1952 152
rect 1956 148 1957 152
rect 1951 147 1957 148
rect 1968 123 1972 152
rect 1975 148 1976 152
rect 1980 148 1981 152
rect 1975 147 1981 148
rect 2176 143 2180 152
rect 2175 142 2181 143
rect 2175 138 2176 142
rect 2180 138 2181 142
rect 2175 137 2181 138
rect 1863 122 1869 123
rect 1863 118 1864 122
rect 1868 118 1869 122
rect 1863 117 1869 118
rect 1967 122 1973 123
rect 1967 118 1968 122
rect 1972 118 1973 122
rect 1967 117 1973 118
rect 2969 92 3033 198
rect 1847 81 1853 82
rect 1847 77 1848 81
rect 1852 77 1853 81
rect 1847 76 1853 77
rect 1695 72 1701 73
rect 1695 68 1696 72
rect 1700 68 1701 72
rect 1695 67 1701 68
rect 1671 62 1677 63
rect 1671 58 1672 62
rect 1676 58 1677 62
rect 1671 57 1677 58
rect 1503 12 1509 13
rect 1503 8 1504 12
rect 1508 8 1509 12
rect 1503 7 1509 8
rect 369 -32 433 -2
rect 1672 1 1676 57
rect 1696 37 1700 67
rect 1712 23 1716 46
rect 1840 33 1844 48
rect 1848 38 1852 76
rect 2015 62 2021 63
rect 2015 58 2016 62
rect 2020 58 2021 62
rect 2969 58 3033 88
rect 3059 1212 3123 1342
rect 3059 1102 3123 1208
rect 3059 992 3123 1098
rect 3059 882 3123 988
rect 3059 772 3123 878
rect 3059 662 3123 768
rect 3059 552 3123 658
rect 3059 442 3123 548
rect 3059 332 3123 438
rect 3059 222 3123 328
rect 3059 112 3123 218
rect 2015 57 2021 58
rect 1839 32 1845 33
rect 1839 28 1840 32
rect 1844 28 1845 32
rect 1839 27 1845 28
rect 1711 22 1717 23
rect 1711 18 1712 22
rect 1716 18 1717 22
rect 1711 17 1717 18
rect 1864 13 1868 46
rect 1952 43 1956 45
rect 1976 43 1980 51
rect 2016 48 2020 57
rect 1951 42 1957 43
rect 1975 42 1981 43
rect 1951 38 1952 42
rect 1956 38 1957 42
rect 1951 37 1957 38
rect 1968 13 1972 42
rect 1975 38 1976 42
rect 1980 38 1981 42
rect 1975 37 1981 38
rect 2176 33 2180 42
rect 2175 32 2181 33
rect 2175 28 2176 32
rect 2180 28 2181 32
rect 2175 27 2181 28
rect 1863 12 1869 13
rect 1863 8 1864 12
rect 1868 8 1869 12
rect 1863 7 1869 8
rect 1967 12 1973 13
rect 1967 8 1968 12
rect 1972 8 1973 12
rect 1967 7 1973 8
rect 3059 2 3123 108
rect 3059 -32 3123 -2
<< m3contact >>
rect 559 2457 563 2461
rect 512 2347 516 2351
rect 504 2237 508 2241
rect 497 2127 501 2131
rect 490 2017 494 2021
rect 483 1907 487 1911
rect 476 1797 480 1801
rect 469 1687 473 1691
rect 462 1577 466 1581
rect 552 1218 556 1222
rect 544 1198 548 1202
rect 559 958 563 962
rect 566 2447 570 2451
rect 662 2737 666 2741
rect 662 2457 666 2461
rect 614 2447 618 2451
rect 590 2347 594 2351
rect 590 2237 594 2241
rect 590 2127 594 2131
rect 590 2017 594 2021
rect 590 1907 594 1911
rect 590 1797 594 1801
rect 846 2457 850 2461
rect 798 2447 802 2451
rect 1030 2457 1034 2461
rect 982 2447 986 2451
rect 774 2347 778 2351
rect 958 2347 962 2351
rect 774 2237 778 2241
rect 774 2127 778 2131
rect 774 2017 778 2021
rect 774 1907 778 1911
rect 774 1797 778 1801
rect 590 1687 594 1691
rect 774 1687 778 1691
rect 590 1577 594 1581
rect 774 1577 778 1581
rect 636 1481 640 1485
rect 566 948 570 952
rect 616 1218 620 1222
rect 643 1471 647 1475
rect 650 1460 654 1464
rect 650 1258 654 1262
rect 657 1450 661 1454
rect 643 1148 647 1152
rect 657 1178 661 1182
rect 665 1440 669 1444
rect 665 1168 669 1172
rect 665 1158 669 1162
rect 672 1430 676 1434
rect 672 1278 676 1282
rect 672 1128 676 1132
rect 680 1420 684 1424
rect 680 1068 684 1072
rect 688 1410 692 1414
rect 657 1058 661 1062
rect 958 2237 962 2241
rect 958 2127 962 2131
rect 958 2017 962 2021
rect 958 1907 962 1911
rect 958 1797 962 1801
rect 958 1687 962 1691
rect 958 1577 962 1581
rect 1070 1541 1074 1545
rect 1094 1481 1098 1485
rect 1086 1471 1090 1475
rect 1078 1460 1082 1464
rect 934 1450 938 1454
rect 926 1440 930 1444
rect 918 1430 922 1434
rect 910 1420 914 1424
rect 902 1410 906 1414
rect 704 1399 708 1403
rect 894 1399 898 1403
rect 688 1048 692 1052
rect 696 1388 700 1392
rect 636 1038 640 1042
rect 664 958 668 962
rect 616 948 620 952
rect 704 1018 708 1022
rect 712 1378 716 1382
rect 696 938 700 942
rect 512 848 516 852
rect 592 848 596 852
rect 560 828 564 832
rect 520 808 524 812
rect 704 828 708 832
rect 552 798 556 802
rect 504 738 508 742
rect 592 738 596 742
rect 560 718 564 722
rect 520 698 524 702
rect 704 718 708 722
rect 552 688 556 692
rect 497 628 501 632
rect 592 628 596 632
rect 560 608 564 612
rect 520 588 524 592
rect 704 608 708 612
rect 720 1368 724 1372
rect 552 578 556 582
rect 490 518 494 522
rect 592 518 596 522
rect 560 498 564 502
rect 520 478 524 482
rect 704 498 708 502
rect 728 1358 732 1362
rect 552 468 556 472
rect 483 408 487 412
rect 592 408 596 412
rect 560 388 564 392
rect 520 368 524 372
rect 704 388 708 392
rect 736 1348 740 1352
rect 552 358 556 362
rect 476 298 480 302
rect 592 298 596 302
rect 560 278 564 282
rect 520 258 524 262
rect 704 278 708 282
rect 744 1338 748 1342
rect 552 248 556 252
rect 469 188 473 192
rect 592 188 596 192
rect 560 168 564 172
rect 520 148 524 152
rect 704 168 708 172
rect 752 1328 756 1332
rect 552 138 556 142
rect 462 78 466 82
rect 592 78 596 82
rect 560 58 564 62
rect 520 38 524 42
rect 704 58 708 62
rect 792 1318 796 1322
rect 768 1258 772 1262
rect 768 1148 772 1152
rect 768 1038 772 1042
rect 960 1308 964 1312
rect 800 1278 804 1282
rect 800 1168 804 1172
rect 800 1058 804 1062
rect 816 958 820 962
rect 1552 958 1556 962
rect 768 948 772 952
rect 1504 948 1508 952
rect 872 938 876 942
rect 1656 868 1660 872
rect 1670 868 1674 872
rect 768 848 772 852
rect 1592 838 1596 842
rect 1616 838 1620 842
rect 912 818 916 822
rect 904 808 908 812
rect 1656 828 1660 832
rect 1672 828 1676 832
rect 1504 778 1508 782
rect 1624 759 1628 763
rect 768 738 772 742
rect 1592 728 1596 732
rect 1616 728 1620 732
rect 912 708 916 712
rect 904 698 908 702
rect 1760 958 1764 962
rect 1712 948 1716 952
rect 1912 958 1916 962
rect 1864 948 1868 952
rect 2080 1198 2084 1202
rect 2144 958 2148 962
rect 2096 948 2100 952
rect 1848 847 1852 851
rect 1696 838 1700 842
rect 2016 828 2020 832
rect 1840 798 1844 802
rect 1712 788 1716 792
rect 1952 808 1956 812
rect 1976 808 1980 812
rect 2176 798 2180 802
rect 1864 778 1868 782
rect 1968 778 1972 782
rect 1688 759 1692 763
rect 1624 718 1628 722
rect 1656 718 1660 722
rect 1848 737 1852 741
rect 1696 728 1700 732
rect 1672 718 1676 722
rect 1504 668 1508 672
rect 768 628 772 632
rect 1592 618 1596 622
rect 1616 618 1620 622
rect 912 598 916 602
rect 904 588 908 592
rect 2016 718 2020 722
rect 1840 688 1844 692
rect 1712 678 1716 682
rect 1952 698 1956 702
rect 1976 698 1980 702
rect 2176 688 2180 692
rect 1864 668 1868 672
rect 1968 668 1972 672
rect 1656 608 1660 612
rect 1848 627 1852 631
rect 1696 618 1700 622
rect 1672 608 1676 612
rect 1504 558 1508 562
rect 768 518 772 522
rect 1592 508 1596 512
rect 1616 508 1620 512
rect 912 488 916 492
rect 904 478 908 482
rect 2016 608 2020 612
rect 1840 578 1844 582
rect 1712 568 1716 572
rect 1952 588 1956 592
rect 1976 588 1980 592
rect 2176 578 2180 582
rect 1864 558 1868 562
rect 1968 558 1972 562
rect 1656 498 1660 502
rect 1848 517 1852 521
rect 1696 508 1700 512
rect 1672 498 1676 502
rect 1504 448 1508 452
rect 768 408 772 412
rect 1592 398 1596 402
rect 1616 398 1620 402
rect 912 378 916 382
rect 904 368 908 372
rect 2016 498 2020 502
rect 1840 468 1844 472
rect 1712 458 1716 462
rect 1952 478 1956 482
rect 1976 478 1980 482
rect 2176 468 2180 472
rect 1864 448 1868 452
rect 1968 448 1972 452
rect 1656 388 1660 392
rect 1848 407 1852 411
rect 1696 398 1700 402
rect 1672 388 1676 392
rect 1504 338 1508 342
rect 768 298 772 302
rect 1592 288 1596 292
rect 1616 288 1620 292
rect 912 268 916 272
rect 904 258 908 262
rect 2016 388 2020 392
rect 1840 358 1844 362
rect 1712 348 1716 352
rect 1952 368 1956 372
rect 1976 368 1980 372
rect 2176 358 2180 362
rect 1864 338 1868 342
rect 1968 338 1972 342
rect 1656 278 1660 282
rect 1848 297 1852 301
rect 1696 288 1700 292
rect 1672 278 1676 282
rect 1504 228 1508 232
rect 768 188 772 192
rect 1592 178 1596 182
rect 1616 178 1620 182
rect 912 158 916 162
rect 904 148 908 152
rect 2016 278 2020 282
rect 1840 248 1844 252
rect 1712 238 1716 242
rect 1952 258 1956 262
rect 1976 258 1980 262
rect 2176 248 2180 252
rect 1864 228 1868 232
rect 1968 228 1972 232
rect 1656 168 1660 172
rect 1504 118 1508 122
rect 768 78 772 82
rect 1592 68 1596 72
rect 1616 68 1620 72
rect 912 48 916 52
rect 904 38 908 42
rect 552 28 556 32
rect 1656 58 1660 62
rect 1848 187 1852 191
rect 1696 178 1700 182
rect 1672 168 1676 172
rect 2016 168 2020 172
rect 1840 138 1844 142
rect 1712 128 1716 132
rect 1952 148 1956 152
rect 1976 148 1980 152
rect 2176 138 2180 142
rect 1864 118 1868 122
rect 1968 118 1972 122
rect 1848 77 1852 81
rect 1696 68 1700 72
rect 1672 58 1676 62
rect 1504 8 1508 12
rect 2016 58 2020 62
rect 1840 28 1844 32
rect 1712 18 1716 22
rect 1952 38 1956 42
rect 1976 38 1980 42
rect 2176 28 2180 32
rect 1864 8 1868 12
rect 1968 8 1972 12
<< metal3 >>
rect 565 2741 667 2742
rect 565 2737 662 2741
rect 666 2737 667 2741
rect 565 2736 667 2737
rect 558 2461 1096 2462
rect 558 2457 559 2461
rect 563 2457 662 2461
rect 666 2457 846 2461
rect 850 2457 1030 2461
rect 1034 2457 1096 2461
rect 558 2456 1096 2457
rect 565 2451 1096 2452
rect 565 2447 566 2451
rect 570 2447 614 2451
rect 618 2447 798 2451
rect 802 2447 982 2451
rect 986 2447 1096 2451
rect 565 2446 1096 2447
rect 511 2351 1096 2352
rect 511 2347 512 2351
rect 516 2347 590 2351
rect 594 2347 774 2351
rect 778 2347 958 2351
rect 962 2347 1096 2351
rect 511 2346 1096 2347
rect 503 2241 1096 2242
rect 503 2237 504 2241
rect 508 2237 590 2241
rect 594 2237 774 2241
rect 778 2237 958 2241
rect 962 2237 1096 2241
rect 503 2236 1096 2237
rect 496 2131 1096 2132
rect 496 2127 497 2131
rect 501 2127 590 2131
rect 594 2127 774 2131
rect 778 2127 958 2131
rect 962 2127 1096 2131
rect 496 2126 1096 2127
rect 489 2021 1096 2022
rect 489 2017 490 2021
rect 494 2017 590 2021
rect 594 2017 774 2021
rect 778 2017 958 2021
rect 962 2017 1096 2021
rect 489 2016 1096 2017
rect 482 1911 1096 1912
rect 482 1907 483 1911
rect 487 1907 590 1911
rect 594 1907 774 1911
rect 778 1907 958 1911
rect 962 1907 1096 1911
rect 482 1906 1096 1907
rect 475 1801 1096 1802
rect 475 1797 476 1801
rect 480 1797 590 1801
rect 594 1797 774 1801
rect 778 1797 958 1801
rect 962 1797 1096 1801
rect 475 1796 1096 1797
rect 468 1691 1096 1692
rect 468 1687 469 1691
rect 473 1687 590 1691
rect 594 1687 774 1691
rect 778 1687 958 1691
rect 962 1687 1096 1691
rect 468 1686 1096 1687
rect 461 1581 1096 1582
rect 461 1577 462 1581
rect 466 1577 590 1581
rect 594 1577 774 1581
rect 778 1577 958 1581
rect 962 1577 1096 1581
rect 461 1576 1096 1577
rect 1069 1545 1206 1546
rect 1069 1541 1070 1545
rect 1074 1541 1206 1545
rect 1069 1540 1206 1541
rect 635 1485 1099 1486
rect 635 1481 636 1485
rect 640 1481 1094 1485
rect 1098 1481 1099 1485
rect 635 1480 1099 1481
rect 642 1475 1091 1476
rect 642 1471 643 1475
rect 647 1471 1086 1475
rect 1090 1471 1091 1475
rect 642 1470 1091 1471
rect 649 1464 1083 1465
rect 649 1460 650 1464
rect 654 1460 1078 1464
rect 1082 1460 1083 1464
rect 649 1459 1083 1460
rect 656 1454 939 1455
rect 656 1450 657 1454
rect 661 1450 934 1454
rect 938 1450 939 1454
rect 656 1449 939 1450
rect 664 1444 931 1445
rect 664 1440 665 1444
rect 669 1440 926 1444
rect 930 1440 931 1444
rect 664 1439 931 1440
rect 671 1434 923 1435
rect 671 1430 672 1434
rect 676 1430 918 1434
rect 922 1430 923 1434
rect 671 1429 923 1430
rect 679 1424 915 1425
rect 679 1420 680 1424
rect 684 1420 910 1424
rect 914 1420 915 1424
rect 679 1419 915 1420
rect 687 1414 907 1415
rect 687 1410 688 1414
rect 692 1410 902 1414
rect 906 1410 907 1414
rect 687 1409 907 1410
rect 703 1403 899 1404
rect 703 1399 704 1403
rect 708 1399 894 1403
rect 898 1399 899 1403
rect 703 1398 899 1399
rect 695 1392 786 1393
rect 695 1388 696 1392
rect 700 1388 786 1392
rect 695 1387 786 1388
rect 711 1382 802 1383
rect 711 1378 712 1382
rect 716 1378 802 1382
rect 711 1377 802 1378
rect 719 1372 810 1373
rect 719 1368 720 1372
rect 724 1368 810 1372
rect 719 1367 810 1368
rect 727 1362 824 1363
rect 727 1358 728 1362
rect 732 1358 824 1362
rect 727 1357 824 1358
rect 735 1352 832 1353
rect 735 1348 736 1352
rect 740 1348 832 1352
rect 735 1347 832 1348
rect 743 1342 840 1343
rect 743 1338 744 1342
rect 748 1338 840 1342
rect 743 1337 840 1338
rect 751 1332 956 1333
rect 751 1328 752 1332
rect 756 1328 956 1332
rect 751 1327 956 1328
rect 791 1322 996 1323
rect 791 1318 792 1322
rect 796 1318 996 1322
rect 791 1317 996 1318
rect 959 1312 996 1313
rect 959 1308 960 1312
rect 964 1308 996 1312
rect 959 1307 996 1308
rect 671 1282 805 1283
rect 671 1278 672 1282
rect 676 1278 800 1282
rect 804 1278 805 1282
rect 671 1277 805 1278
rect 649 1262 773 1263
rect 649 1258 650 1262
rect 654 1258 768 1262
rect 772 1258 773 1262
rect 649 1257 773 1258
rect 551 1222 956 1223
rect 551 1218 552 1222
rect 556 1218 616 1222
rect 620 1218 956 1222
rect 551 1217 956 1218
rect 543 1202 2085 1203
rect 543 1198 544 1202
rect 548 1198 2080 1202
rect 2084 1198 2085 1202
rect 543 1197 2085 1198
rect 656 1182 892 1183
rect 656 1178 657 1182
rect 661 1178 892 1182
rect 656 1177 892 1178
rect 664 1172 805 1173
rect 664 1168 665 1172
rect 669 1168 800 1172
rect 804 1168 805 1172
rect 664 1167 805 1168
rect 664 1162 860 1163
rect 664 1158 665 1162
rect 669 1158 860 1162
rect 664 1157 860 1158
rect 642 1152 773 1153
rect 642 1148 643 1152
rect 647 1148 768 1152
rect 772 1148 773 1152
rect 642 1147 773 1148
rect 671 1132 828 1133
rect 671 1128 672 1132
rect 676 1128 828 1132
rect 671 1127 828 1128
rect 679 1072 892 1073
rect 679 1068 680 1072
rect 684 1068 892 1072
rect 679 1067 892 1068
rect 656 1062 805 1063
rect 656 1058 657 1062
rect 661 1058 800 1062
rect 804 1058 805 1062
rect 656 1057 805 1058
rect 687 1052 860 1053
rect 687 1048 688 1052
rect 692 1048 860 1052
rect 687 1047 860 1048
rect 635 1042 773 1043
rect 635 1038 636 1042
rect 640 1038 768 1042
rect 772 1038 773 1042
rect 635 1037 773 1038
rect 703 1022 828 1023
rect 703 1018 704 1022
rect 708 1018 828 1022
rect 703 1017 828 1018
rect 558 962 2149 963
rect 558 958 559 962
rect 563 958 664 962
rect 668 958 816 962
rect 820 958 1552 962
rect 1556 958 1760 962
rect 1764 958 1912 962
rect 1916 958 2144 962
rect 2148 958 2149 962
rect 558 957 2149 958
rect 565 952 2101 953
rect 565 948 566 952
rect 570 948 616 952
rect 620 948 768 952
rect 772 948 1504 952
rect 1508 948 1712 952
rect 1716 948 1864 952
rect 1868 948 2096 952
rect 2100 948 2101 952
rect 565 947 2101 948
rect 695 942 877 943
rect 695 938 696 942
rect 700 938 872 942
rect 876 938 877 942
rect 695 937 877 938
rect 1655 872 1675 873
rect 1655 868 1656 872
rect 1660 868 1670 872
rect 1674 868 1675 872
rect 1655 867 1675 868
rect 502 852 773 853
rect 502 848 512 852
rect 516 848 592 852
rect 596 848 768 852
rect 772 848 773 852
rect 502 847 773 848
rect 1847 851 2186 853
rect 1847 847 1848 851
rect 1852 847 2186 851
rect 1847 846 1853 847
rect 503 842 1621 843
rect 503 838 1592 842
rect 1596 838 1616 842
rect 1620 838 1621 842
rect 503 837 1621 838
rect 1695 842 2186 843
rect 1695 838 1696 842
rect 1700 838 2186 842
rect 1695 837 2186 838
rect 503 832 565 833
rect 503 828 560 832
rect 564 828 565 832
rect 503 827 565 828
rect 703 832 1661 833
rect 703 828 704 832
rect 708 828 1656 832
rect 1660 828 1661 832
rect 703 827 1661 828
rect 1671 832 2021 833
rect 1671 828 1672 832
rect 1676 828 2016 832
rect 2020 828 2021 832
rect 1671 827 2021 828
rect 911 822 925 823
rect 911 818 912 822
rect 916 818 925 822
rect 911 817 925 818
rect 519 812 1981 813
rect 519 808 520 812
rect 524 808 904 812
rect 908 808 1952 812
rect 1956 808 1976 812
rect 1980 808 1981 812
rect 519 807 1981 808
rect 551 802 2181 803
rect 551 798 552 802
rect 556 798 1840 802
rect 1844 798 2176 802
rect 2180 798 2181 802
rect 551 797 2181 798
rect 1487 792 1717 793
rect 1487 788 1712 792
rect 1716 788 1717 792
rect 1487 787 1717 788
rect 1487 782 1509 783
rect 1487 778 1504 782
rect 1508 778 1509 782
rect 1487 777 1509 778
rect 1863 782 2186 783
rect 1863 778 1864 782
rect 1868 778 1968 782
rect 1972 778 2186 782
rect 1863 777 2186 778
rect 1623 763 1693 764
rect 1623 759 1624 763
rect 1628 759 1688 763
rect 1692 759 1693 763
rect 1623 758 1693 759
rect 349 742 773 743
rect 349 738 504 742
rect 508 738 592 742
rect 596 738 768 742
rect 772 738 773 742
rect 349 737 773 738
rect 1847 741 2186 743
rect 1847 737 1848 741
rect 1852 737 2186 741
rect 1847 736 1853 737
rect 503 732 1621 733
rect 503 728 1592 732
rect 1596 728 1616 732
rect 1620 728 1621 732
rect 503 727 1621 728
rect 1695 732 2186 733
rect 1695 728 1696 732
rect 1700 728 2186 732
rect 1695 727 2186 728
rect 503 722 565 723
rect 503 718 560 722
rect 564 718 565 722
rect 503 717 565 718
rect 703 722 1661 723
rect 703 718 704 722
rect 708 718 1624 722
rect 1628 718 1656 722
rect 1660 718 1661 722
rect 703 717 1661 718
rect 1671 722 2021 723
rect 1671 718 1672 722
rect 1676 718 2016 722
rect 2020 718 2021 722
rect 1671 717 2021 718
rect 911 712 925 713
rect 911 708 912 712
rect 916 708 925 712
rect 911 707 925 708
rect 519 702 1981 703
rect 519 698 520 702
rect 524 698 904 702
rect 908 698 1952 702
rect 1956 698 1976 702
rect 1980 698 1981 702
rect 519 697 1981 698
rect 551 692 2181 693
rect 551 688 552 692
rect 556 688 1840 692
rect 1844 688 2176 692
rect 2180 688 2181 692
rect 551 687 2181 688
rect 1487 682 1717 683
rect 1487 678 1712 682
rect 1716 678 1717 682
rect 1487 677 1717 678
rect 1487 672 1509 673
rect 1487 668 1504 672
rect 1508 668 1509 672
rect 1487 667 1509 668
rect 1863 672 2186 673
rect 1863 668 1864 672
rect 1868 668 1968 672
rect 1972 668 2186 672
rect 1863 667 2186 668
rect 342 632 773 633
rect 342 628 497 632
rect 501 628 592 632
rect 596 628 768 632
rect 772 628 773 632
rect 342 627 773 628
rect 1847 631 2186 633
rect 1847 627 1848 631
rect 1852 627 2186 631
rect 1847 626 1853 627
rect 503 622 1621 623
rect 503 618 1592 622
rect 1596 618 1616 622
rect 1620 618 1621 622
rect 503 617 1621 618
rect 1695 622 2186 623
rect 1695 618 1696 622
rect 1700 618 2186 622
rect 1695 617 2186 618
rect 503 612 565 613
rect 503 608 560 612
rect 564 608 565 612
rect 503 607 565 608
rect 703 612 1661 613
rect 703 608 704 612
rect 708 608 1656 612
rect 1660 608 1661 612
rect 703 607 1661 608
rect 1671 612 2021 613
rect 1671 608 1672 612
rect 1676 608 2016 612
rect 2020 608 2021 612
rect 1671 607 2021 608
rect 911 602 925 603
rect 911 598 912 602
rect 916 598 925 602
rect 911 597 925 598
rect 519 592 1981 593
rect 519 588 520 592
rect 524 588 904 592
rect 908 588 1952 592
rect 1956 588 1976 592
rect 1980 588 1981 592
rect 519 587 1981 588
rect 551 582 2181 583
rect 551 578 552 582
rect 556 578 1840 582
rect 1844 578 2176 582
rect 2180 578 2181 582
rect 551 577 2181 578
rect 1487 572 1717 573
rect 1487 568 1712 572
rect 1716 568 1717 572
rect 1487 567 1717 568
rect 1487 562 1509 563
rect 1487 558 1504 562
rect 1508 558 1509 562
rect 1487 557 1509 558
rect 1863 562 2186 563
rect 1863 558 1864 562
rect 1868 558 1968 562
rect 1972 558 2186 562
rect 1863 557 2186 558
rect 343 522 773 523
rect 343 518 490 522
rect 494 518 592 522
rect 596 518 768 522
rect 772 518 773 522
rect 343 517 773 518
rect 1847 521 2186 523
rect 1847 517 1848 521
rect 1852 517 2186 521
rect 1847 516 1853 517
rect 503 512 1621 513
rect 503 508 1592 512
rect 1596 508 1616 512
rect 1620 508 1621 512
rect 503 507 1621 508
rect 1695 512 2186 513
rect 1695 508 1696 512
rect 1700 508 2186 512
rect 1695 507 2186 508
rect 503 502 565 503
rect 503 498 560 502
rect 564 498 565 502
rect 503 497 565 498
rect 703 502 1661 503
rect 703 498 704 502
rect 708 498 1656 502
rect 1660 498 1661 502
rect 703 497 1661 498
rect 1671 502 2021 503
rect 1671 498 1672 502
rect 1676 498 2016 502
rect 2020 498 2021 502
rect 1671 497 2021 498
rect 911 492 925 493
rect 911 488 912 492
rect 916 488 925 492
rect 911 487 925 488
rect 519 482 1981 483
rect 519 478 520 482
rect 524 478 904 482
rect 908 478 1952 482
rect 1956 478 1976 482
rect 1980 478 1981 482
rect 519 477 1981 478
rect 551 472 2181 473
rect 551 468 552 472
rect 556 468 1840 472
rect 1844 468 2176 472
rect 2180 468 2181 472
rect 551 467 2181 468
rect 1487 462 1717 463
rect 1487 458 1712 462
rect 1716 458 1717 462
rect 1487 457 1717 458
rect 1487 452 1509 453
rect 1487 448 1504 452
rect 1508 448 1509 452
rect 1487 447 1509 448
rect 1863 452 2186 453
rect 1863 448 1864 452
rect 1868 448 1968 452
rect 1972 448 2186 452
rect 1863 447 2186 448
rect 342 412 773 413
rect 342 408 483 412
rect 487 408 592 412
rect 596 408 768 412
rect 772 408 773 412
rect 342 407 773 408
rect 1847 411 2186 413
rect 1847 407 1848 411
rect 1852 407 2186 411
rect 1847 406 1853 407
rect 503 402 1621 403
rect 503 398 1592 402
rect 1596 398 1616 402
rect 1620 398 1621 402
rect 503 397 1621 398
rect 1695 402 2186 403
rect 1695 398 1696 402
rect 1700 398 2186 402
rect 1695 397 2186 398
rect 503 392 565 393
rect 503 388 560 392
rect 564 388 565 392
rect 503 387 565 388
rect 703 392 1661 393
rect 703 388 704 392
rect 708 388 1656 392
rect 1660 388 1661 392
rect 703 387 1661 388
rect 1671 392 2021 393
rect 1671 388 1672 392
rect 1676 388 2016 392
rect 2020 388 2021 392
rect 1671 387 2021 388
rect 911 382 925 383
rect 911 378 912 382
rect 916 378 925 382
rect 911 377 925 378
rect 519 372 1981 373
rect 519 368 520 372
rect 524 368 904 372
rect 908 368 1952 372
rect 1956 368 1976 372
rect 1980 368 1981 372
rect 519 367 1981 368
rect 551 362 2181 363
rect 551 358 552 362
rect 556 358 1840 362
rect 1844 358 2176 362
rect 2180 358 2181 362
rect 551 357 2181 358
rect 1487 352 1717 353
rect 1487 348 1712 352
rect 1716 348 1717 352
rect 1487 347 1717 348
rect 1487 342 1509 343
rect 1487 338 1504 342
rect 1508 338 1509 342
rect 1487 337 1509 338
rect 1863 342 2186 343
rect 1863 338 1864 342
rect 1868 338 1968 342
rect 1972 338 2186 342
rect 1863 337 2186 338
rect 340 302 773 303
rect 340 298 476 302
rect 480 298 592 302
rect 596 298 768 302
rect 772 298 773 302
rect 340 297 773 298
rect 1847 301 2186 303
rect 1847 297 1848 301
rect 1852 297 2186 301
rect 1847 296 1853 297
rect 503 292 1621 293
rect 503 288 1592 292
rect 1596 288 1616 292
rect 1620 288 1621 292
rect 503 287 1621 288
rect 1695 292 2186 293
rect 1695 288 1696 292
rect 1700 288 2186 292
rect 1695 287 2186 288
rect 503 282 565 283
rect 503 278 560 282
rect 564 278 565 282
rect 503 277 565 278
rect 703 282 1661 283
rect 703 278 704 282
rect 708 278 1656 282
rect 1660 278 1661 282
rect 703 277 1661 278
rect 1671 282 2021 283
rect 1671 278 1672 282
rect 1676 278 2016 282
rect 2020 278 2021 282
rect 1671 277 2021 278
rect 911 272 925 273
rect 911 268 912 272
rect 916 268 925 272
rect 911 267 925 268
rect 519 262 1981 263
rect 519 258 520 262
rect 524 258 904 262
rect 908 258 1952 262
rect 1956 258 1976 262
rect 1980 258 1981 262
rect 519 257 1981 258
rect 551 252 2181 253
rect 551 248 552 252
rect 556 248 1840 252
rect 1844 248 2176 252
rect 2180 248 2181 252
rect 551 247 2181 248
rect 1487 242 1717 243
rect 1487 238 1712 242
rect 1716 238 1717 242
rect 1487 237 1717 238
rect 1487 232 1509 233
rect 1487 228 1504 232
rect 1508 228 1509 232
rect 1487 227 1509 228
rect 1863 232 2186 233
rect 1863 228 1864 232
rect 1868 228 1968 232
rect 1972 228 2186 232
rect 1863 227 2186 228
rect 339 192 773 193
rect 339 188 469 192
rect 473 188 592 192
rect 596 188 768 192
rect 772 188 773 192
rect 339 187 773 188
rect 1847 191 2186 193
rect 1847 187 1848 191
rect 1852 187 2186 191
rect 1847 186 1853 187
rect 503 182 1621 183
rect 503 178 1592 182
rect 1596 178 1616 182
rect 1620 178 1621 182
rect 503 177 1621 178
rect 1695 182 2186 183
rect 1695 178 1696 182
rect 1700 178 2186 182
rect 1695 177 2186 178
rect 503 172 565 173
rect 503 168 560 172
rect 564 168 565 172
rect 503 167 565 168
rect 703 172 1661 173
rect 703 168 704 172
rect 708 168 1656 172
rect 1660 168 1661 172
rect 703 167 1661 168
rect 1671 172 2021 173
rect 1671 168 1672 172
rect 1676 168 2016 172
rect 2020 168 2021 172
rect 1671 167 2021 168
rect 911 162 925 163
rect 911 158 912 162
rect 916 158 925 162
rect 911 157 925 158
rect 519 152 1981 153
rect 519 148 520 152
rect 524 148 904 152
rect 908 148 1952 152
rect 1956 148 1976 152
rect 1980 148 1981 152
rect 519 147 1981 148
rect 551 142 2181 143
rect 551 138 552 142
rect 556 138 1840 142
rect 1844 138 2176 142
rect 2180 138 2181 142
rect 551 137 2181 138
rect 1487 132 1717 133
rect 1487 128 1712 132
rect 1716 128 1717 132
rect 1487 127 1717 128
rect 1487 122 1509 123
rect 1487 118 1504 122
rect 1508 118 1509 122
rect 1487 117 1509 118
rect 1863 122 2186 123
rect 1863 118 1864 122
rect 1868 118 1968 122
rect 1972 118 2186 122
rect 1863 117 2186 118
rect 339 82 773 83
rect 339 78 462 82
rect 466 78 592 82
rect 596 78 768 82
rect 772 78 773 82
rect 339 77 773 78
rect 1847 81 2186 83
rect 1847 77 1848 81
rect 1852 77 2186 81
rect 1847 76 1853 77
rect 503 72 1621 73
rect 503 68 1592 72
rect 1596 68 1616 72
rect 1620 68 1621 72
rect 503 67 1621 68
rect 1695 72 2186 73
rect 1695 68 1696 72
rect 1700 68 2186 72
rect 1695 67 2186 68
rect 503 62 565 63
rect 503 58 560 62
rect 564 58 565 62
rect 503 57 565 58
rect 703 62 1661 63
rect 703 58 704 62
rect 708 58 1656 62
rect 1660 58 1661 62
rect 703 57 1661 58
rect 1671 62 2021 63
rect 1671 58 1672 62
rect 1676 58 2016 62
rect 2020 58 2021 62
rect 1671 57 2021 58
rect 911 52 925 53
rect 911 48 912 52
rect 916 48 925 52
rect 911 47 925 48
rect 519 42 1981 43
rect 519 38 520 42
rect 524 38 904 42
rect 908 38 1952 42
rect 1956 38 1976 42
rect 1980 38 1981 42
rect 519 37 1981 38
rect 551 32 2181 33
rect 551 28 552 32
rect 556 28 1840 32
rect 1844 28 2176 32
rect 2180 28 2181 32
rect 551 27 2181 28
rect 1487 22 1717 23
rect 1487 18 1712 22
rect 1716 18 1717 22
rect 1487 17 1717 18
rect 1487 12 1509 13
rect 1487 8 1504 12
rect 1508 8 1509 12
rect 1487 7 1509 8
rect 1863 12 2186 13
rect 1863 8 1864 12
rect 1868 8 1968 12
rect 1972 8 2186 12
rect 1863 7 2186 8
use flopen_1x_8  flopen_1x_8_0
timestamp 1493660808
transform 1 0 574 0 1 1499
box -6 -4 138 976
use flopen_1x_8  flopen_1x_8_1
timestamp 1493660808
transform 1 0 758 0 1 1499
box -6 -4 138 976
use flopen_1x_8  flopen_1x_8_2
timestamp 1493660808
transform 1 0 942 0 1 1499
box -6 -4 138 976
use mux2_c_1x  mux2_c_1x_0
timestamp 1492902181
transform 1 0 760 0 1 1210
box -6 -4 66 96
use mux2_c_1x  mux2_c_1x_1
timestamp 1492902181
transform 1 0 760 0 1 1100
box -6 -4 66 96
use mux2_c_1x  mux2_c_1x_2
timestamp 1492902181
transform 1 0 760 0 1 990
box -6 -4 66 96
use mux2_1x_8  mux2_1x_8_0
timestamp 1484532969
transform 1 0 520 0 1 0
box -6 -4 50 976
use flopen_1x_8  flopen_1x_8_3
timestamp 1493660808
transform 1 0 576 0 1 0
box -6 -4 138 976
use flop_1x_8  flop_1x_8_0
timestamp 1484532171
transform 1 0 761 0 1 0
box -7 -4 105 976
use mux2_1x_8  mux2_1x_8_1
timestamp 1484532969
transform 1 0 872 0 1 0
box -6 -4 50 976
use flop_1x_8  flop_1x_8_1
timestamp 1484532171
transform 1 0 1497 0 1 0
box -7 -4 105 976
use mux4_1x_8  mux4_1x_8_0
timestamp 1484532969
transform 1 0 1600 0 1 0
box -6 -4 106 976
use flop_1x_8  flop_1x_8_2
timestamp 1484532171
transform 1 0 1705 0 1 0
box -7 -4 105 976
use mux2_1x_8  mux2_1x_8_2
timestamp 1484532969
transform 1 0 1808 0 1 0
box -6 -4 50 976
use flop_1x_8  flop_1x_8_3
timestamp 1484532171
transform 1 0 1857 0 1 0
box -7 -4 105 976
use mux3_1x_8  mux3_1x_8_0
timestamp 1484532969
transform 1 0 1960 0 1 0
box -6 -4 82 976
use flopenr_1x_8  flopenr_1x_8_0
timestamp 1484532171
transform 1 0 2040 0 1 0
box -6 -4 147 976
use alt_alu  alt_alu_0
timestamp 1493063752
transform 1 0 2217 0 1 -4
box -33 0 377 986
use shifter  shifter_0
timestamp 1492982022
transform 1 0 2761 0 1 -4
box -172 0 192 1648
use regramarray_dp  regramarray_dp_0
timestamp 1488938149
transform 1 0 920 0 1 0
box -102 -5 578 1306
<< labels >>
rlabel metal2 2218 1309 2218 1309 1 zero
rlabel metal2 2050 1309 2050 1309 1 pcen
rlabel metal2 1994 1310 1994 1310 1 pcsrc_1_
rlabel metal2 1962 1309 1962 1309 1 pcsrc_0
rlabel metal2 1809 1309 1809 1309 1 alusrca
rlabel metal2 1633 1310 1633 1310 1 alusrcb_1_
rlabel metal2 1601 1310 1601 1310 1 alusrcb_0_
rlabel m3contact 961 1310 961 1310 1 regwrite
rlabel metal2 3090 1316 3090 1316 1 Gnd!
rlabel metal2 3000 1327 3000 1327 1 Vdd!
rlabel m2contact 2751 1640 2755 1644 5 op8
rlabel m2contact 2808 1640 2812 1644 5 op7
rlabel metal2 2273 1310 2273 1310 1 op6
rlabel metal2 2281 1310 2281 1310 1 op5
rlabel metal2 2313 1310 2313 1310 1 op4
rlabel metal2 2329 1310 2329 1310 1 op3
rlabel metal2 2346 1310 2346 1310 1 op2
rlabel metal2 2465 1310 2465 1310 1 op0
rlabel metal2 2505 1310 2505 1310 1 op1
rlabel metal3 2182 850 2182 850 1 a7
rlabel metal3 2182 840 2182 840 1 b7
rlabel metal3 2181 780 2181 780 1 result7
rlabel metal3 2181 740 2181 740 1 a6
rlabel metal3 2181 730 2181 730 1 b6
rlabel metal3 2181 670 2181 670 1 result6
rlabel metal3 2181 630 2181 630 1 a5
rlabel metal3 2181 620 2181 620 1 b5
rlabel metal3 2180 560 2180 560 1 result5
rlabel metal3 2180 520 2180 520 1 a4
rlabel metal3 2180 510 2180 510 1 b4
rlabel metal3 2179 450 2179 450 1 result4
rlabel metal3 2179 410 2179 410 1 a3
rlabel metal3 2179 400 2179 400 1 b3
rlabel metal3 2181 340 2181 340 1 result3
rlabel metal3 2180 300 2180 300 1 a2
rlabel metal3 2180 290 2180 290 1 b2
rlabel metal3 2180 230 2180 230 1 result2
rlabel metal3 2181 190 2181 190 1 a1
rlabel metal3 2181 180 2181 180 1 b1
rlabel metal3 2181 120 2181 120 1 result1
rlabel metal3 2181 80 2181 80 1 a0
rlabel metal3 2181 70 2181 70 1 b0
rlabel metal3 2181 10 2181 10 1 result0
rlabel metal2 586 1310 586 1310 1 irwrite_0_
rlabel metal2 698 1310 698 1310 1 memtoreg
rlabel metal2 714 1309 714 1309 1 funct_5_
rlabel metal2 722 1310 722 1310 1 funct_4_
rlabel metal2 730 1309 730 1309 1 funct_3_
rlabel metal2 738 1311 738 1311 1 funct_2_
rlabel metal2 746 1308 746 1308 1 funct_1_
rlabel metal2 753 1309 753 1309 1 funct_0_
rlabel metal2 522 1310 522 1310 1 iord
rlabel metal3 505 60 505 60 1 adr0
rlabel metal3 505 70 505 70 1 writedata0
rlabel metal3 506 80 506 80 1 memdata0
rlabel metal3 505 170 505 170 1 adr1
rlabel metal3 505 180 505 180 1 writedata1
rlabel metal3 506 190 506 190 1 memdata1
rlabel metal3 506 280 506 280 1 adr2
rlabel metal3 506 290 506 290 1 writedata2
rlabel metal3 507 300 507 300 1 memdata2
rlabel metal3 506 390 506 390 1 adr3
rlabel metal3 507 400 507 400 1 writedata3
rlabel metal3 506 409 506 409 1 memdata3
rlabel metal3 506 500 506 500 1 adr4
rlabel metal3 506 510 506 510 1 writedata4
rlabel metal3 506 519 506 519 1 memdata4
rlabel metal3 505 610 505 610 1 adr5
rlabel metal3 505 619 505 619 1 writedata5
rlabel metal3 506 630 506 630 1 memdata5
rlabel metal3 506 721 506 721 1 adr6
rlabel metal3 505 729 505 729 1 writedata6
rlabel m3contact 505 739 505 739 1 memdata6
rlabel metal3 507 831 507 831 1 adr7
rlabel metal3 507 839 507 839 1 writedata7
rlabel metal3 507 850 507 850 1 memdata7
rlabel metal2 794 1309 794 1309 1 regdst
rlabel metal3 568 2739 568 2739 1 ph1
rlabel metal2 584 2809 584 2809 1 irwrite_3_
rlabel metal2 712 2808 712 2808 1 op_5_
rlabel metal2 720 2809 720 2809 1 op_4_
rlabel metal2 728 2808 728 2808 1 op_3_
rlabel metal2 736 2810 736 2810 1 op_2_
rlabel metal2 744 2807 744 2807 1 op_1_
rlabel metal2 752 2809 752 2809 1 op_0_
rlabel metal2 768 2809 768 2809 1 irwrite_2_
rlabel metal2 952 2809 952 2809 1 irwrite_1_
rlabel metal2 554 1309 554 1309 1 ph2
rlabel metal2 546 1308 546 1308 1 reset
rlabel metal2 397 1326 397 1326 1 Gnd!
rlabel metal2 309 1327 309 1327 1 Vdd!
rlabel metal2 2807 1310 2811 1314 1 s2
rlabel metal2 2871 1092 2875 1096 1 s1
rlabel metal2 2919 984 2923 988 1 s0
rlabel metal2 1690 1034 1690 1034 1 shamt0
rlabel metal2 1672 1034 1672 1034 1 shamt1
rlabel metal3 1203 1543 1203 1543 1 shamt2
<< end >>
