magic
tech scmos
timestamp 1492456146
<< metal1 >>
rect -66 1142 -50 1146
rect -66 1032 -58 1036
rect -46 930 -42 934
rect -66 922 -50 926
rect -2 922 6 926
rect -54 820 -38 824
rect -66 812 -58 816
rect -2 812 6 816
rect -46 710 -42 714
rect -66 702 -50 706
rect -2 702 6 706
rect -54 600 -38 604
rect -66 592 -58 596
rect -2 592 6 596
rect -46 490 -42 494
rect -66 482 -50 486
rect -2 482 6 486
rect -54 380 -38 384
rect -66 372 -58 376
rect -2 372 6 376
rect -46 270 -42 274
rect -66 262 -50 266
rect -2 262 6 266
rect -54 160 -38 164
rect -2 152 6 156
rect -52 90 -43 98
rect -46 50 -42 54
rect -53 0 -44 8
<< m2contact >>
rect -50 1142 -46 1146
rect -58 1032 -54 1036
rect -50 930 -46 934
rect -50 922 -46 926
rect 6 922 10 926
rect -58 820 -54 824
rect -58 812 -54 816
rect 6 812 10 816
rect -50 710 -46 714
rect -50 702 -46 706
rect 6 702 10 706
rect -58 600 -54 604
rect -58 592 -54 596
rect 6 592 10 596
rect -50 490 -46 494
rect -50 482 -46 486
rect 6 482 10 486
rect -58 380 -54 384
rect -58 372 -54 376
rect 6 372 10 376
rect -50 270 -46 274
rect -50 262 -46 266
rect 6 262 10 266
rect -58 160 -54 164
rect 6 152 10 156
rect -50 50 -46 54
<< metal2 >>
rect -66 915 -62 926
rect -58 824 -54 1032
rect -50 934 -46 1142
rect -66 805 -62 816
rect -66 695 -62 706
rect -58 604 -54 812
rect -50 714 -46 922
rect -10 915 -6 932
rect -10 805 -6 822
rect 6 820 10 922
rect 38 816 42 822
rect -66 585 -62 596
rect -66 475 -62 486
rect -58 384 -54 592
rect -50 494 -46 702
rect -10 695 -6 712
rect 6 710 10 812
rect 38 706 42 712
rect -10 585 -6 602
rect 6 600 10 702
rect 38 596 42 602
rect -66 365 -62 376
rect -66 255 -62 266
rect -58 164 -54 372
rect -50 274 -46 482
rect -10 475 -6 492
rect 6 490 10 592
rect 38 486 42 492
rect -10 365 -6 382
rect 6 380 10 482
rect 38 376 42 382
rect -66 145 -62 156
rect -50 54 -46 262
rect -10 255 -6 272
rect 6 270 10 372
rect 38 266 42 272
rect -10 145 -6 162
rect 6 160 10 262
rect 38 156 42 162
rect -66 35 -62 46
rect -10 35 -6 52
rect 6 50 10 152
rect 38 46 42 52
<< m3contact >>
rect -66 911 -62 915
rect -66 801 -62 805
rect -66 691 -62 695
rect -10 911 -6 915
rect -10 801 -6 805
rect 6 812 10 816
rect 38 812 42 816
rect -66 581 -62 585
rect -66 471 -62 475
rect -10 691 -6 695
rect 6 702 10 706
rect 38 702 42 706
rect -10 581 -6 585
rect 6 592 10 596
rect 38 592 42 596
rect -66 361 -62 365
rect -66 251 -62 255
rect -10 471 -6 475
rect 6 482 10 486
rect 38 482 42 486
rect -10 361 -6 365
rect 6 372 10 376
rect 38 372 42 376
rect -66 141 -62 145
rect -10 251 -6 255
rect 6 262 10 266
rect 38 262 42 266
rect -10 141 -6 145
rect 6 152 10 156
rect 38 152 42 156
rect -66 31 -62 35
rect -2 42 2 46
rect 38 42 42 46
rect -10 31 -6 35
<< metal3 >>
rect -67 915 -5 916
rect -67 911 -66 915
rect -62 911 -10 915
rect -6 911 -5 915
rect -67 910 -5 911
rect 5 816 43 817
rect 5 812 6 816
rect 10 812 38 816
rect 42 812 43 816
rect 5 811 43 812
rect -67 805 -5 806
rect -67 801 -66 805
rect -62 801 -10 805
rect -6 801 -5 805
rect -67 800 -5 801
rect 5 706 43 707
rect 5 702 6 706
rect 10 702 38 706
rect 42 702 43 706
rect 5 701 43 702
rect -67 695 -5 696
rect -67 691 -66 695
rect -62 691 -10 695
rect -6 691 -5 695
rect -67 690 -5 691
rect 5 596 43 597
rect 5 592 6 596
rect 10 592 38 596
rect 42 592 43 596
rect 5 591 43 592
rect -67 585 -5 586
rect -67 581 -66 585
rect -62 581 -10 585
rect -6 581 -5 585
rect -67 580 -5 581
rect 5 486 43 487
rect 5 482 6 486
rect 10 482 38 486
rect 42 482 43 486
rect 5 481 43 482
rect -67 475 -5 476
rect -67 471 -66 475
rect -62 471 -10 475
rect -6 471 -5 475
rect -67 470 -5 471
rect 5 376 43 377
rect 5 372 6 376
rect 10 372 38 376
rect 42 372 43 376
rect 5 371 43 372
rect -67 365 -5 366
rect -67 361 -66 365
rect -62 361 -10 365
rect -6 361 -5 365
rect -67 360 -5 361
rect 5 266 43 267
rect 5 262 6 266
rect 10 262 38 266
rect 42 262 43 266
rect 5 261 43 262
rect -67 255 -5 256
rect -67 251 -66 255
rect -62 251 -10 255
rect -6 251 -5 255
rect -67 250 -5 251
rect 5 156 43 157
rect 5 152 6 156
rect 10 152 38 156
rect 42 152 43 156
rect 5 151 43 152
rect -67 145 -5 146
rect -67 141 -66 145
rect -62 141 -10 145
rect -6 141 -5 145
rect -67 140 -5 141
rect -3 46 43 47
rect -3 42 -2 46
rect 2 42 38 46
rect 42 42 43 46
rect -3 41 43 42
rect -67 35 -5 36
rect -67 31 -66 35
rect -62 31 -10 35
rect -6 31 -5 35
rect -67 30 -5 31
use mux2_dp_1x  mux2_dp_1x_6
timestamp 1484435125
transform 1 0 -106 0 1 1104
box -6 -4 50 96
use mux2_dp_1x  mux2_dp_1x_5
timestamp 1484435125
transform 1 0 -106 0 1 994
box -6 -4 50 96
use mux2_dp_1x  mux2_dp_1x_4
timestamp 1484435125
transform 1 0 -106 0 1 884
box -6 -4 50 96
use mux2_dp_1x  mux2_dp_1x_3
timestamp 1484435125
transform 1 0 -42 0 1 884
box -6 -4 50 96
use mux2_dp_1x  mux2_dp_1x_2
array 1 1 56 1 8 110
timestamp 1484435125
transform 1 0 -106 0 1 4
box -6 -4 50 96
use mux2_dp_1x  mux2_dp_1x_1
array 1 1 56 1 8 110
timestamp 1484435125
transform 1 0 -42 0 1 4
box -6 -4 50 96
use mux2_dp_1x  mux2_dp_1x_0
array 1 1 56 1 8 110
timestamp 1484435125
transform 1 0 6 0 1 4
box -6 -4 50 96
<< end >>
