magic
tech scmos
timestamp 1488310061
<< nwell >>
rect -9 48 26 105
<< ntransistor >>
rect 7 6 9 26
<< ptransistor >>
rect 7 54 9 94
<< ndiffusion >>
rect 2 25 7 26
rect 6 6 7 25
rect 9 25 14 26
rect 9 6 10 25
<< pdiffusion >>
rect 2 93 7 94
rect 6 54 7 93
rect 9 93 14 94
rect 9 54 10 93
<< ndcontact >>
rect 2 6 6 25
rect 10 6 14 25
<< pdcontact >>
rect 2 54 6 93
rect 10 54 14 93
<< psubstratepcontact >>
rect -2 -2 2 2
<< nsubstratencontact >>
rect -2 98 2 102
<< polysilicon >>
rect 7 94 9 96
rect 7 33 9 54
rect 6 29 9 33
rect 7 26 9 29
rect 7 4 9 6
<< polycontact >>
rect 2 29 6 33
<< metal1 >>
rect -2 102 18 103
rect 2 98 18 102
rect -2 97 18 98
rect 2 93 6 97
rect 10 93 14 94
rect 2 33 6 37
rect 2 25 6 26
rect 10 25 14 54
rect 2 3 6 6
rect -2 2 18 3
rect 2 -2 18 2
rect -2 -3 18 -2
<< labels >>
flabel metal1 4 100 4 100 4 FreeSans 26 0 0 0 vdd
flabel metal1 4 0 4 0 4 FreeSans 26 0 0 0 gnd
flabel metal1 12 45 12 45 4 FreeSans 26 0 0 0 Y
flabel metal1 4 35 4 35 4 FreeSans 26 0 0 0 A
<< end >>
