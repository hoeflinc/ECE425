magic
tech scmos
timestamp 1488306862
<< m2contact >>
rect -2 -2 2 2
<< end >>
