.subckt inv a y N=4 P=8
M1 y a gnd gnd NMOS W='N' L=2 
+ AS='N*5' PS='2*N+10' AD='N*5' PD='2*N+10'
M2 y a vdddriver vdddriver PMOS W='P' L=2
+ AS='P*5' PS='2*P+10' AD='P*5' PD='2*P+10'
.ends
