magic
tech scmos
timestamp 1488310061
<< m2contact >>
rect -2 -2 2 2
<< end >>
