magic
tech scmos
timestamp 1493661823
<< metal2 >>
rect -33 1621 -27 1622
rect -33 1617 -32 1621
rect -28 1617 -27 1621
rect -33 1616 -27 1617
rect -41 1602 -35 1603
rect -41 1598 -40 1602
rect -36 1598 -35 1602
rect -41 1597 -35 1598
rect -243 1278 -179 1343
rect -123 1308 -119 1312
rect -40 1308 -36 1597
rect -32 1308 -28 1616
rect -25 1572 -19 1573
rect -25 1568 -24 1572
rect -20 1568 -19 1572
rect -25 1567 -19 1568
rect -24 1308 -20 1567
rect 0 1308 4 1312
rect 56 1308 60 1312
rect 184 1308 188 1312
rect 192 1308 196 1312
rect 200 1308 204 1312
rect 208 1308 212 1312
rect 216 1308 220 1312
rect 224 1308 228 1312
rect 240 1308 244 1312
rect 424 1308 428 1312
rect 584 1308 588 1312
rect 696 1308 700 1312
rect 728 1308 732 1312
rect 736 1308 740 1312
rect 744 1308 748 1312
rect 752 1308 756 1312
rect 792 1308 796 1312
rect 960 1308 964 1312
rect 1600 1308 1604 1312
rect 1632 1308 1636 1312
rect 1808 1308 1812 1312
rect 1960 1308 1964 1312
rect 1992 1308 1996 1312
rect 2048 1308 2052 1312
rect 2216 1308 2220 1312
rect 2240 1308 2244 1312
rect 2480 1308 2484 1312
rect 2512 1308 2516 1312
rect 2634 1278 2698 1862
rect 2724 1278 2788 1863
<< m3contact >>
rect -32 1617 -28 1621
rect -40 1598 -36 1602
rect -24 1568 -20 1572
rect -12 1428 -8 1432
rect -16 848 -12 852
rect -16 838 -12 842
rect -16 828 -12 832
rect -16 738 -12 742
rect -16 728 -12 732
rect -16 718 -12 722
rect -16 628 -12 632
rect -16 618 -12 622
rect -16 608 -12 612
rect -16 518 -12 522
rect -16 508 -12 512
rect -16 498 -12 502
rect -16 408 -12 412
rect -16 398 -12 402
rect -16 388 -12 392
rect -16 298 -12 302
rect -16 288 -12 292
rect -16 278 -12 282
rect -16 188 -12 192
rect -16 178 -12 182
rect -16 168 -12 172
rect -16 78 -12 82
rect -16 68 -12 72
rect -16 58 -12 62
<< metal3 >>
rect -63 1621 -27 1622
rect -63 1617 -32 1621
rect -28 1617 -27 1621
rect -63 1616 -27 1617
rect -63 1602 -35 1603
rect -63 1598 -40 1602
rect -36 1598 -35 1602
rect -63 1597 -35 1598
rect -63 1572 -19 1573
rect -63 1568 -24 1572
rect -20 1568 -19 1572
rect -63 1567 -19 1568
use controller  controller_0
timestamp 1492976468
transform 1 0 0 0 1 1450
box -243 -172 2788 368
use datapath  datapath_0
timestamp 1493661823
transform 1 0 0 0 1 0
box -243 -32 2788 1343
<< labels >>
rlabel metal3 -62 1598 -58 1602 1 reset
rlabel metal3 -62 1568 -58 1572 1 ph2
rlabel metal3 -62 1617 -58 1621 1 ph1
rlabel m3contact -12 1428 -8 1432 1 memwrite
rlabel m3contact -16 848 -12 852 1 memdata7
rlabel m3contact -16 838 -12 842 1 writedata7
rlabel m3contact -16 828 -12 832 1 adr7
rlabel m3contact -16 738 -12 742 1 memdata6
rlabel m3contact -16 728 -12 732 1 writedata6
rlabel m3contact -16 718 -12 722 1 adr6
rlabel m3contact -16 628 -12 632 1 memdata5
rlabel m3contact -16 618 -12 622 1 writedata5
rlabel m3contact -16 608 -12 612 1 adr5
rlabel m3contact -16 518 -12 522 1 memdata4
rlabel m3contact -16 508 -12 512 1 writedata4
rlabel m3contact -16 498 -12 502 1 adr4
rlabel m3contact -16 408 -12 412 1 memdata3
rlabel m3contact -16 398 -12 402 1 writedata3
rlabel m3contact -16 388 -12 392 1 adr3
rlabel m3contact -16 298 -12 302 1 memdata2
rlabel m3contact -16 288 -12 292 1 writedata2
rlabel m3contact -16 278 -12 282 1 adr2
rlabel m3contact -16 188 -12 192 1 memdata1
rlabel m3contact -16 178 -12 182 1 writedata1
rlabel m3contact -16 168 -12 172 1 adr1
rlabel m3contact -16 78 -12 82 1 memdata0
rlabel m3contact -16 68 -12 72 1 writedata0
rlabel m3contact -16 58 -12 62 1 adr0
<< end >>
