magic
tech scmos
timestamp 1493953340
<< metal1 >>
rect -98 1296 510 1304
rect -98 1206 510 1214
rect -98 1186 518 1194
rect -98 1096 518 1104
rect -98 1076 518 1084
rect -98 986 518 994
rect 22 966 534 974
rect 38 876 550 884
rect 70 856 509 864
rect -2 766 509 774
rect 70 746 509 754
rect -2 656 509 664
rect 70 636 509 644
rect -2 546 509 554
rect 70 526 509 534
rect -2 436 509 444
rect 70 416 509 424
rect -2 326 509 334
rect 70 306 509 314
rect -2 216 509 224
rect 70 196 509 204
rect -2 106 509 114
rect 70 86 509 94
rect -2 3 77 4
rect 142 3 509 4
rect -2 -4 509 3
rect 70 -5 149 -4
<< metal2 >>
rect -9 1292 -3 1293
rect -9 1288 -8 1292
rect -4 1288 -3 1292
rect -9 1287 -3 1288
rect 71 1292 77 1293
rect 71 1288 72 1292
rect 76 1288 77 1292
rect 71 1287 77 1288
rect 215 1292 221 1293
rect 215 1288 216 1292
rect 220 1288 221 1292
rect 215 1287 221 1288
rect 359 1292 365 1293
rect 359 1288 360 1292
rect 364 1288 365 1292
rect 359 1287 365 1288
rect 503 1292 509 1293
rect 503 1288 504 1292
rect 508 1288 509 1292
rect 503 1287 509 1288
rect -25 1282 -19 1283
rect -25 1278 -24 1282
rect -20 1278 -19 1282
rect -25 1277 -19 1278
rect -41 1272 -35 1273
rect -41 1268 -40 1272
rect -36 1268 -35 1272
rect -41 1267 -35 1268
rect -57 1262 -51 1263
rect -57 1258 -56 1262
rect -52 1258 -51 1262
rect -57 1257 -51 1258
rect -96 1248 -92 1252
rect -88 1233 -84 1251
rect -72 1243 -68 1251
rect -64 1248 -60 1252
rect -56 1249 -52 1257
rect -40 1249 -36 1267
rect -32 1248 -28 1252
rect -24 1249 -20 1277
rect -8 1249 -4 1287
rect -1 1282 5 1283
rect -1 1278 0 1282
rect 4 1278 5 1282
rect -1 1277 5 1278
rect 0 1264 4 1277
rect 7 1262 13 1263
rect 7 1258 8 1262
rect 12 1258 13 1262
rect 7 1257 13 1258
rect 8 1255 12 1257
rect -73 1242 -67 1243
rect -73 1238 -72 1242
rect -68 1238 -67 1242
rect -73 1237 -67 1238
rect 16 1233 20 1257
rect -89 1232 -83 1233
rect -89 1228 -88 1232
rect -84 1228 -83 1232
rect -89 1227 -83 1228
rect 15 1232 21 1233
rect 15 1228 16 1232
rect 20 1228 21 1232
rect 15 1227 21 1228
rect 32 1223 36 1257
rect 40 1253 44 1266
rect 72 1264 76 1287
rect 143 1282 149 1283
rect 143 1278 144 1282
rect 148 1278 149 1282
rect 143 1277 149 1278
rect 79 1262 85 1263
rect 79 1258 80 1262
rect 84 1258 85 1262
rect 79 1257 85 1258
rect 80 1255 84 1257
rect 39 1252 45 1253
rect 39 1248 40 1252
rect 44 1248 45 1252
rect 39 1247 45 1248
rect 88 1233 92 1257
rect 87 1232 93 1233
rect 87 1228 88 1232
rect 92 1228 93 1232
rect 87 1227 93 1228
rect 104 1223 108 1257
rect 112 1253 116 1266
rect 144 1264 148 1277
rect 151 1272 157 1273
rect 151 1268 152 1272
rect 156 1268 157 1272
rect 151 1267 157 1268
rect 152 1255 156 1267
rect 111 1252 117 1253
rect 111 1248 112 1252
rect 116 1248 117 1252
rect 111 1247 117 1248
rect 160 1233 164 1257
rect 159 1232 165 1233
rect 159 1228 160 1232
rect 164 1228 165 1232
rect 159 1227 165 1228
rect 176 1223 180 1257
rect 184 1253 188 1266
rect 216 1264 220 1287
rect 287 1282 293 1283
rect 287 1278 288 1282
rect 292 1278 293 1282
rect 287 1277 293 1278
rect 223 1272 229 1273
rect 223 1268 224 1272
rect 228 1268 229 1272
rect 223 1267 229 1268
rect 224 1255 228 1267
rect 183 1252 189 1253
rect 183 1248 184 1252
rect 188 1248 189 1252
rect 183 1247 189 1248
rect 232 1233 236 1257
rect 231 1232 237 1233
rect 231 1228 232 1232
rect 236 1228 237 1232
rect 231 1227 237 1228
rect 248 1223 252 1257
rect 256 1253 260 1266
rect 288 1264 292 1277
rect 295 1262 301 1263
rect 295 1258 296 1262
rect 300 1258 301 1262
rect 295 1257 301 1258
rect 296 1255 300 1257
rect 255 1252 261 1253
rect 255 1248 256 1252
rect 260 1248 261 1252
rect 255 1247 261 1248
rect 304 1243 308 1257
rect 303 1242 309 1243
rect 303 1238 304 1242
rect 308 1238 309 1242
rect 303 1237 309 1238
rect 320 1223 324 1257
rect 328 1253 332 1266
rect 360 1264 364 1287
rect 431 1282 437 1283
rect 431 1278 432 1282
rect 436 1278 437 1282
rect 431 1277 437 1278
rect 367 1262 373 1263
rect 367 1258 368 1262
rect 372 1258 373 1262
rect 367 1257 373 1258
rect 368 1255 372 1257
rect 327 1252 333 1253
rect 327 1248 328 1252
rect 332 1248 333 1252
rect 327 1247 333 1248
rect 376 1243 380 1257
rect 375 1242 381 1243
rect 375 1238 376 1242
rect 380 1238 381 1242
rect 375 1237 381 1238
rect 392 1223 396 1257
rect 400 1253 404 1266
rect 432 1264 436 1277
rect 439 1272 445 1273
rect 439 1268 440 1272
rect 444 1268 445 1272
rect 439 1267 445 1268
rect 440 1255 444 1267
rect 399 1252 405 1253
rect 399 1248 400 1252
rect 404 1248 405 1252
rect 399 1247 405 1248
rect 448 1243 452 1257
rect 447 1242 453 1243
rect 447 1238 448 1242
rect 452 1238 453 1242
rect 447 1237 453 1238
rect 464 1223 468 1257
rect 472 1253 476 1266
rect 504 1264 508 1287
rect 511 1272 517 1273
rect 511 1268 512 1272
rect 516 1268 517 1272
rect 511 1267 517 1268
rect 512 1255 516 1267
rect 471 1252 477 1253
rect 471 1248 472 1252
rect 476 1248 477 1252
rect 471 1247 477 1248
rect 520 1243 524 1257
rect 519 1242 525 1243
rect 519 1238 520 1242
rect 524 1238 525 1242
rect 519 1237 525 1238
rect 536 1223 540 1257
rect 544 1253 548 1266
rect 543 1252 549 1253
rect 543 1248 544 1252
rect 548 1248 549 1252
rect 543 1247 549 1248
rect 31 1222 37 1223
rect 31 1218 32 1222
rect 36 1218 37 1222
rect 31 1217 37 1218
rect 103 1222 109 1223
rect 103 1218 104 1222
rect 108 1218 109 1222
rect 103 1217 109 1218
rect 175 1222 181 1223
rect 175 1218 176 1222
rect 180 1218 181 1222
rect 175 1217 181 1218
rect 247 1222 253 1223
rect 247 1218 248 1222
rect 252 1218 253 1222
rect 247 1217 253 1218
rect 319 1222 325 1223
rect 319 1218 320 1222
rect 324 1218 325 1222
rect 319 1217 325 1218
rect 391 1222 397 1223
rect 391 1218 392 1222
rect 396 1218 397 1222
rect 391 1217 397 1218
rect 463 1222 469 1223
rect 463 1218 464 1222
rect 468 1218 469 1222
rect 463 1217 469 1218
rect 535 1222 541 1223
rect 535 1218 536 1222
rect 540 1218 541 1222
rect 535 1217 541 1218
rect -33 1182 -27 1183
rect -33 1178 -32 1182
rect -28 1178 -27 1182
rect -33 1177 -27 1178
rect -9 1182 -3 1183
rect -9 1178 -8 1182
rect -4 1178 -3 1182
rect -9 1177 -3 1178
rect 79 1182 85 1183
rect 79 1178 80 1182
rect 84 1178 85 1182
rect 79 1177 85 1178
rect 223 1182 229 1183
rect 223 1178 224 1182
rect 228 1178 229 1182
rect 223 1177 229 1178
rect 367 1182 373 1183
rect 367 1178 368 1182
rect 372 1178 373 1182
rect 367 1177 373 1178
rect 511 1182 517 1183
rect 511 1178 512 1182
rect 516 1178 517 1182
rect 511 1177 517 1178
rect -65 1162 -59 1163
rect -65 1158 -64 1162
rect -60 1158 -59 1162
rect -65 1157 -59 1158
rect -41 1162 -35 1163
rect -41 1158 -40 1162
rect -36 1158 -35 1162
rect -41 1157 -35 1158
rect -96 1133 -92 1141
rect -97 1132 -91 1133
rect -97 1128 -96 1132
rect -92 1128 -91 1132
rect -97 1127 -91 1128
rect -88 1123 -84 1141
rect -72 1133 -68 1141
rect -64 1139 -60 1157
rect -57 1152 -51 1153
rect -57 1148 -56 1152
rect -52 1148 -51 1152
rect -57 1147 -51 1148
rect -56 1139 -52 1147
rect -40 1139 -36 1157
rect -32 1139 -28 1177
rect -25 1172 -19 1173
rect -25 1168 -24 1172
rect -20 1168 -19 1172
rect -25 1167 -19 1168
rect -24 1139 -20 1167
rect -8 1139 -4 1177
rect 7 1172 13 1173
rect 7 1168 8 1172
rect 12 1168 13 1172
rect 7 1167 13 1168
rect 8 1144 12 1167
rect 15 1152 21 1153
rect 15 1148 16 1152
rect 20 1148 21 1152
rect 15 1147 21 1148
rect 16 1144 20 1147
rect -73 1132 -67 1133
rect -73 1128 -72 1132
rect -68 1128 -67 1132
rect -73 1127 -67 1128
rect 24 1123 28 1146
rect 80 1144 84 1177
rect 151 1172 157 1173
rect 151 1168 152 1172
rect 156 1168 157 1172
rect 151 1167 157 1168
rect 87 1152 93 1153
rect 87 1148 88 1152
rect 92 1148 93 1152
rect 87 1147 93 1148
rect 88 1144 92 1147
rect 96 1123 100 1146
rect 152 1144 156 1167
rect 159 1162 165 1163
rect 159 1158 160 1162
rect 164 1158 165 1162
rect 159 1157 165 1158
rect 160 1144 164 1157
rect 168 1123 172 1146
rect 224 1144 228 1177
rect 295 1172 301 1173
rect 295 1168 296 1172
rect 300 1168 301 1172
rect 295 1167 301 1168
rect 231 1162 237 1163
rect 231 1158 232 1162
rect 236 1158 237 1162
rect 231 1157 237 1158
rect 232 1144 236 1157
rect 240 1123 244 1146
rect 296 1144 300 1167
rect 303 1152 309 1153
rect 303 1148 304 1152
rect 308 1148 309 1152
rect 303 1147 309 1148
rect 304 1144 308 1147
rect 312 1133 316 1146
rect 368 1144 372 1177
rect 439 1172 445 1173
rect 439 1168 440 1172
rect 444 1168 445 1172
rect 439 1167 445 1168
rect 375 1152 381 1153
rect 375 1148 376 1152
rect 380 1148 381 1152
rect 375 1147 381 1148
rect 376 1144 380 1147
rect 384 1133 388 1146
rect 440 1144 444 1167
rect 447 1162 453 1163
rect 447 1158 448 1162
rect 452 1158 453 1162
rect 447 1157 453 1158
rect 448 1144 452 1157
rect 456 1133 460 1146
rect 512 1144 516 1177
rect 519 1162 525 1163
rect 519 1158 520 1162
rect 524 1158 525 1162
rect 519 1157 525 1158
rect 520 1144 524 1157
rect 528 1133 532 1146
rect 311 1132 317 1133
rect 311 1128 312 1132
rect 316 1128 317 1132
rect 311 1127 317 1128
rect 383 1132 389 1133
rect 383 1128 384 1132
rect 388 1128 389 1132
rect 383 1127 389 1128
rect 455 1132 461 1133
rect 455 1128 456 1132
rect 460 1128 461 1132
rect 455 1127 461 1128
rect 527 1132 533 1133
rect 527 1128 528 1132
rect 532 1128 533 1132
rect 527 1127 533 1128
rect -89 1122 -83 1123
rect -89 1118 -88 1122
rect -84 1118 -83 1122
rect -89 1117 -83 1118
rect 23 1122 29 1123
rect 23 1118 24 1122
rect 28 1118 29 1122
rect 23 1117 29 1118
rect 95 1122 101 1123
rect 95 1118 96 1122
rect 100 1118 101 1122
rect 95 1117 101 1118
rect 167 1122 173 1123
rect 167 1118 168 1122
rect 172 1118 173 1122
rect 167 1117 173 1118
rect 239 1122 245 1123
rect 239 1118 240 1122
rect 244 1118 245 1122
rect 239 1117 245 1118
rect -33 1072 -27 1073
rect -33 1068 -32 1072
rect -28 1068 -27 1072
rect -33 1067 -27 1068
rect -9 1072 -3 1073
rect -9 1068 -8 1072
rect -4 1068 -3 1072
rect -9 1067 -3 1068
rect 79 1072 85 1073
rect 79 1068 80 1072
rect 84 1068 85 1072
rect 79 1067 85 1068
rect 223 1072 229 1073
rect 223 1068 224 1072
rect 228 1068 229 1072
rect 223 1067 229 1068
rect 367 1072 373 1073
rect 367 1068 368 1072
rect 372 1068 373 1072
rect 367 1067 373 1068
rect 511 1072 517 1073
rect 511 1068 512 1072
rect 516 1068 517 1072
rect 511 1067 517 1068
rect -65 1052 -59 1053
rect -65 1048 -64 1052
rect -60 1048 -59 1052
rect -65 1047 -59 1048
rect -41 1052 -35 1053
rect -41 1048 -40 1052
rect -36 1048 -35 1052
rect -41 1047 -35 1048
rect -96 1023 -92 1031
rect -97 1022 -91 1023
rect -97 1018 -96 1022
rect -92 1018 -91 1022
rect -97 1017 -91 1018
rect -88 1013 -84 1031
rect -72 1023 -68 1031
rect -64 1029 -60 1047
rect -57 1042 -51 1043
rect -57 1038 -56 1042
rect -52 1038 -51 1042
rect -57 1037 -51 1038
rect -56 1029 -52 1037
rect -40 1029 -36 1047
rect -32 1029 -28 1067
rect -25 1062 -19 1063
rect -25 1058 -24 1062
rect -20 1058 -19 1062
rect -25 1057 -19 1058
rect -24 1029 -20 1057
rect -8 1029 -4 1067
rect 7 1062 13 1063
rect 7 1058 8 1062
rect 12 1058 13 1062
rect 7 1057 13 1058
rect 8 1034 12 1057
rect 15 1042 21 1043
rect 15 1038 16 1042
rect 20 1038 21 1042
rect 15 1037 21 1038
rect 16 1034 20 1037
rect -73 1022 -67 1023
rect -73 1018 -72 1022
rect -68 1018 -67 1022
rect -73 1017 -67 1018
rect 24 1013 28 1036
rect 80 1034 84 1067
rect 151 1062 157 1063
rect 151 1058 152 1062
rect 156 1058 157 1062
rect 151 1057 157 1058
rect 87 1042 93 1043
rect 87 1038 88 1042
rect 92 1038 93 1042
rect 87 1037 93 1038
rect 88 1034 92 1037
rect 96 1013 100 1036
rect 152 1034 156 1057
rect 159 1052 165 1053
rect 159 1048 160 1052
rect 164 1048 165 1052
rect 159 1047 165 1048
rect 160 1034 164 1047
rect 168 1013 172 1036
rect 224 1034 228 1067
rect 295 1062 301 1063
rect 295 1058 296 1062
rect 300 1058 301 1062
rect 295 1057 301 1058
rect 231 1052 237 1053
rect 231 1048 232 1052
rect 236 1048 237 1052
rect 231 1047 237 1048
rect 232 1034 236 1047
rect 240 1013 244 1036
rect 296 1034 300 1057
rect 303 1042 309 1043
rect 303 1038 304 1042
rect 308 1038 309 1042
rect 303 1037 309 1038
rect 304 1034 308 1037
rect 312 1023 316 1036
rect 368 1034 372 1067
rect 439 1062 445 1063
rect 439 1058 440 1062
rect 444 1058 445 1062
rect 439 1057 445 1058
rect 375 1042 381 1043
rect 375 1038 376 1042
rect 380 1038 381 1042
rect 375 1037 381 1038
rect 376 1034 380 1037
rect 384 1023 388 1036
rect 440 1034 444 1057
rect 447 1052 453 1053
rect 447 1048 448 1052
rect 452 1048 453 1052
rect 447 1047 453 1048
rect 448 1034 452 1047
rect 456 1023 460 1036
rect 512 1034 516 1067
rect 519 1052 525 1053
rect 519 1048 520 1052
rect 524 1048 525 1052
rect 519 1047 525 1048
rect 520 1034 524 1047
rect 528 1023 532 1036
rect 311 1022 317 1023
rect 311 1018 312 1022
rect 316 1018 317 1022
rect 311 1017 317 1018
rect 383 1022 389 1023
rect 383 1018 384 1022
rect 388 1018 389 1022
rect 383 1017 389 1018
rect 455 1022 461 1023
rect 455 1018 456 1022
rect 460 1018 461 1022
rect 455 1017 461 1018
rect 527 1022 533 1023
rect 527 1018 528 1022
rect 532 1018 533 1022
rect 527 1017 533 1018
rect -89 1012 -83 1013
rect -89 1008 -88 1012
rect -84 1008 -83 1012
rect -89 1007 -83 1008
rect 23 1012 29 1013
rect 23 1008 24 1012
rect 28 1008 29 1012
rect 23 1007 29 1008
rect 95 1012 101 1013
rect 95 1008 96 1012
rect 100 1008 101 1012
rect 95 1007 101 1008
rect 167 1012 173 1013
rect 167 1008 168 1012
rect 172 1008 173 1012
rect 167 1007 173 1008
rect 239 1012 245 1013
rect 239 1008 240 1012
rect 244 1008 245 1012
rect 239 1007 245 1008
<< m3contact >>
rect -8 1288 -4 1292
rect 72 1288 76 1292
rect 216 1288 220 1292
rect 360 1288 364 1292
rect 504 1288 508 1292
rect -24 1278 -20 1282
rect -40 1268 -36 1272
rect -56 1258 -52 1262
rect 0 1278 4 1282
rect 8 1258 12 1262
rect -72 1238 -68 1242
rect -88 1228 -84 1232
rect 16 1228 20 1232
rect 144 1278 148 1282
rect 80 1258 84 1262
rect 40 1248 44 1252
rect 88 1228 92 1232
rect 152 1268 156 1272
rect 112 1248 116 1252
rect 160 1228 164 1232
rect 288 1278 292 1282
rect 224 1268 228 1272
rect 184 1248 188 1252
rect 232 1228 236 1232
rect 296 1258 300 1262
rect 256 1248 260 1252
rect 304 1238 308 1242
rect 432 1278 436 1282
rect 368 1258 372 1262
rect 328 1248 332 1252
rect 376 1238 380 1242
rect 440 1268 444 1272
rect 400 1248 404 1252
rect 448 1238 452 1242
rect 512 1268 516 1272
rect 472 1248 476 1252
rect 520 1238 524 1242
rect 544 1248 548 1252
rect 32 1218 36 1222
rect 104 1218 108 1222
rect 176 1218 180 1222
rect 248 1218 252 1222
rect 320 1218 324 1222
rect 392 1218 396 1222
rect 464 1218 468 1222
rect 536 1218 540 1222
rect -32 1178 -28 1182
rect -8 1178 -4 1182
rect 80 1178 84 1182
rect 224 1178 228 1182
rect 368 1178 372 1182
rect 512 1178 516 1182
rect -64 1158 -60 1162
rect -40 1158 -36 1162
rect -96 1128 -92 1132
rect -56 1148 -52 1152
rect -24 1168 -20 1172
rect 8 1168 12 1172
rect 16 1148 20 1152
rect -72 1128 -68 1132
rect 152 1168 156 1172
rect 88 1148 92 1152
rect 160 1158 164 1162
rect 296 1168 300 1172
rect 232 1158 236 1162
rect 304 1148 308 1152
rect 440 1168 444 1172
rect 376 1148 380 1152
rect 448 1158 452 1162
rect 520 1158 524 1162
rect 312 1128 316 1132
rect 384 1128 388 1132
rect 456 1128 460 1132
rect 528 1128 532 1132
rect -88 1118 -84 1122
rect 24 1118 28 1122
rect 96 1118 100 1122
rect 168 1118 172 1122
rect 240 1118 244 1122
rect -32 1068 -28 1072
rect -8 1068 -4 1072
rect 80 1068 84 1072
rect 224 1068 228 1072
rect 368 1068 372 1072
rect 512 1068 516 1072
rect -64 1048 -60 1052
rect -40 1048 -36 1052
rect -96 1018 -92 1022
rect -56 1038 -52 1042
rect -24 1058 -20 1062
rect 8 1058 12 1062
rect 16 1038 20 1042
rect -72 1018 -68 1022
rect 152 1058 156 1062
rect 88 1038 92 1042
rect 160 1048 164 1052
rect 296 1058 300 1062
rect 232 1048 236 1052
rect 304 1038 308 1042
rect 440 1058 444 1062
rect 376 1038 380 1042
rect 448 1048 452 1052
rect 520 1048 524 1052
rect 312 1018 316 1022
rect 384 1018 388 1022
rect 456 1018 460 1022
rect 528 1018 532 1022
rect -88 1008 -84 1012
rect 24 1008 28 1012
rect 96 1008 100 1012
rect 168 1008 172 1012
rect 240 1008 244 1012
<< metal3 >>
rect -9 1292 509 1293
rect -9 1288 -8 1292
rect -4 1288 72 1292
rect 76 1288 216 1292
rect 220 1288 360 1292
rect 364 1288 504 1292
rect 508 1288 509 1292
rect -9 1287 509 1288
rect -25 1282 437 1283
rect -25 1278 -24 1282
rect -20 1278 0 1282
rect 4 1278 144 1282
rect 148 1278 288 1282
rect 292 1278 432 1282
rect 436 1278 437 1282
rect -25 1277 437 1278
rect -41 1272 517 1273
rect -41 1268 -40 1272
rect -36 1268 152 1272
rect 156 1268 224 1272
rect 228 1268 440 1272
rect 444 1268 512 1272
rect 516 1268 517 1272
rect -41 1267 517 1268
rect -57 1262 373 1263
rect -57 1258 -56 1262
rect -52 1258 8 1262
rect 12 1258 80 1262
rect 84 1258 296 1262
rect 300 1258 368 1262
rect 372 1258 373 1262
rect -57 1257 373 1258
rect 39 1252 549 1253
rect 39 1248 40 1252
rect 44 1248 112 1252
rect 116 1248 184 1252
rect 188 1248 256 1252
rect 260 1248 328 1252
rect 332 1248 400 1252
rect 404 1248 472 1252
rect 476 1248 544 1252
rect 548 1248 549 1252
rect 39 1247 549 1248
rect -73 1242 525 1243
rect -73 1238 -72 1242
rect -68 1238 304 1242
rect 308 1238 376 1242
rect 380 1238 448 1242
rect 452 1238 520 1242
rect 524 1238 525 1242
rect -73 1237 525 1238
rect -89 1232 237 1233
rect -89 1228 -88 1232
rect -84 1228 16 1232
rect 20 1228 88 1232
rect 92 1228 160 1232
rect 164 1228 232 1232
rect 236 1228 237 1232
rect -89 1227 237 1228
rect 31 1222 541 1223
rect 31 1218 32 1222
rect 36 1218 104 1222
rect 108 1218 176 1222
rect 180 1218 248 1222
rect 252 1218 320 1222
rect 324 1218 392 1222
rect 396 1218 464 1222
rect 468 1218 536 1222
rect 540 1218 541 1222
rect 31 1217 541 1218
rect -33 1182 -27 1183
rect -33 1178 -32 1182
rect -28 1178 -27 1182
rect -33 1177 -27 1178
rect -9 1182 517 1183
rect -9 1178 -8 1182
rect -4 1178 80 1182
rect 84 1178 224 1182
rect 228 1178 368 1182
rect 372 1178 512 1182
rect 516 1178 517 1182
rect -9 1177 517 1178
rect -25 1172 445 1173
rect -25 1168 -24 1172
rect -20 1168 8 1172
rect 12 1168 152 1172
rect 156 1168 296 1172
rect 300 1168 440 1172
rect 444 1168 445 1172
rect -25 1167 445 1168
rect -65 1162 -59 1163
rect -65 1158 -64 1162
rect -60 1158 -59 1162
rect -65 1157 -59 1158
rect -41 1162 525 1163
rect -41 1158 -40 1162
rect -36 1158 160 1162
rect 164 1158 232 1162
rect 236 1158 448 1162
rect 452 1158 520 1162
rect 524 1158 525 1162
rect -41 1157 525 1158
rect -57 1152 381 1153
rect -57 1148 -56 1152
rect -52 1148 16 1152
rect 20 1148 88 1152
rect 92 1148 304 1152
rect 308 1148 376 1152
rect 380 1148 381 1152
rect -57 1147 381 1148
rect -97 1132 -91 1133
rect -97 1128 -96 1132
rect -92 1128 -91 1132
rect -97 1127 -91 1128
rect -73 1132 533 1133
rect -73 1128 -72 1132
rect -68 1128 312 1132
rect 316 1128 384 1132
rect 388 1128 456 1132
rect 460 1128 528 1132
rect 532 1128 533 1132
rect -73 1127 533 1128
rect -89 1122 245 1123
rect -89 1118 -88 1122
rect -84 1118 24 1122
rect 28 1118 96 1122
rect 100 1118 168 1122
rect 172 1118 240 1122
rect 244 1118 245 1122
rect -89 1117 245 1118
rect -33 1072 -27 1073
rect -33 1068 -32 1072
rect -28 1068 -27 1072
rect -33 1067 -27 1068
rect -9 1072 517 1073
rect -9 1068 -8 1072
rect -4 1068 80 1072
rect 84 1068 224 1072
rect 228 1068 368 1072
rect 372 1068 512 1072
rect 516 1068 517 1072
rect -9 1067 517 1068
rect -25 1062 445 1063
rect -25 1058 -24 1062
rect -20 1058 8 1062
rect 12 1058 152 1062
rect 156 1058 296 1062
rect 300 1058 440 1062
rect 444 1058 445 1062
rect -25 1057 445 1058
rect -65 1052 -59 1053
rect -65 1048 -64 1052
rect -60 1048 -59 1052
rect -65 1047 -59 1048
rect -41 1052 525 1053
rect -41 1048 -40 1052
rect -36 1048 160 1052
rect 164 1048 232 1052
rect 236 1048 448 1052
rect 452 1048 520 1052
rect 524 1048 525 1052
rect -41 1047 525 1048
rect -57 1042 381 1043
rect -57 1038 -56 1042
rect -52 1038 16 1042
rect 20 1038 88 1042
rect 92 1038 304 1042
rect 308 1038 376 1042
rect 380 1038 381 1042
rect -57 1037 381 1038
rect -97 1022 -91 1023
rect -97 1018 -96 1022
rect -92 1018 -91 1022
rect -97 1017 -91 1018
rect -73 1022 533 1023
rect -73 1018 -72 1022
rect -68 1018 312 1022
rect 316 1018 384 1022
rect 388 1018 456 1022
rect 460 1018 528 1022
rect 532 1018 533 1022
rect -73 1017 533 1018
rect -89 1012 245 1013
rect -89 1008 -88 1012
rect -84 1008 24 1012
rect 28 1008 96 1012
rect 100 1008 168 1012
rect 172 1008 240 1012
rect 244 1008 245 1012
rect -89 1007 245 1008
rect -1 817 508 823
rect 39 787 573 793
rect 63 777 573 783
rect -1 707 508 713
rect 39 677 573 683
rect 63 667 573 673
rect -1 597 508 603
rect 39 567 573 573
rect 63 557 573 563
rect -1 487 508 493
rect 39 457 573 463
rect 63 447 573 453
rect -1 377 508 383
rect 39 347 573 353
rect 63 337 573 343
rect -1 267 508 273
rect 39 237 573 243
rect 63 227 573 233
rect -1 157 508 163
rect 39 127 573 133
rect 63 117 573 123
rect -1 47 508 53
rect 39 17 573 23
rect 63 7 573 13
use invbuf_4x  invbuf_4x_0
timestamp 1484532969
transform 1 0 -96 0 1 1210
box -6 -4 34 96
use invbuf_4x  invbuf_4x_1
timestamp 1484532969
transform 1 0 -64 0 1 1210
box -6 -4 34 96
use invbuf_4x  invbuf_4x_2
timestamp 1484532969
transform 1 0 -32 0 1 1210
box -6 -4 34 96
use invbuf_4x  invbuf_4x_3
timestamp 1484532969
transform 1 0 -96 0 1 1100
box -6 -4 34 96
use invbuf_4x  invbuf_4x_4
timestamp 1484532969
transform 1 0 -64 0 1 1100
box -6 -4 34 96
use invbuf_4x  invbuf_4x_5
timestamp 1484532969
transform 1 0 -32 0 1 1100
box -6 -4 34 96
use invbuf_4x  invbuf_4x_6
timestamp 1484532969
transform 1 0 -96 0 1 990
box -6 -4 34 96
use invbuf_4x  invbuf_4x_7
timestamp 1484532969
transform 1 0 -64 0 1 990
box -6 -4 34 96
use invbuf_4x  invbuf_4x_8
timestamp 1484532969
transform 1 0 -32 0 1 990
box -6 -4 34 96
use regramvector0_dp  regramvector0_dp_0
timestamp 1484533619
transform 1 0 0 0 1 0
box -6 -4 74 1306
use regramvector_dp  regramvector_dp_0
timestamp 1484533408
transform 1 0 72 0 1 0
box -6 -4 74 1306
use regramvector_dp  regramvector_dp_1
timestamp 1484533408
transform 1 0 144 0 1 0
box -6 -4 74 1306
use regramvector_dp  regramvector_dp_2
timestamp 1484533408
transform 1 0 216 0 1 0
box -6 -4 74 1306
use regramvector_dp  regramvector_dp_3
timestamp 1484533408
transform 1 0 288 0 1 0
box -6 -4 74 1306
use regramvector_dp  regramvector_dp_4
timestamp 1484533408
transform 1 0 360 0 1 0
box -6 -4 74 1306
use regramvector_dp  regramvector_dp_5
timestamp 1484533408
transform 1 0 432 0 1 0
box -6 -4 74 1306
use regramvector_dp  regramvector_dp_6
timestamp 1484533408
transform 1 0 504 0 1 0
box -6 -4 74 1306
<< labels >>
rlabel metal2 -94 1250 -94 1250 1 wa_2_
rlabel metal2 -62 1250 -62 1250 1 wa_1_
rlabel metal2 -30 1250 -30 1250 1 wa_0_
rlabel m3contact 42 1250 42 1250 1 regwrite
rlabel m3contact -94 1130 -94 1130 1 ra2_2_
rlabel m3contact -94 1020 -94 1020 1 ra1_2_
rlabel m3contact -62 1050 -62 1050 1 ra1_1_
rlabel m3contact -30 1069 -30 1069 1 ra1_0_
rlabel metal3 1 820 1 820 1 w_7_
rlabel metal3 1 710 1 710 1 w_6_
rlabel metal3 1 600 1 600 1 w_5_
rlabel metal3 1 490 1 490 1 w_4_
rlabel metal3 1 380 1 380 1 w_3_
rlabel metal3 1 270 1 270 1 w_2_
rlabel metal3 1 160 1 160 1 w_1_
rlabel metal3 1 50 1 50 1 w_0_
rlabel metal3 570 20 570 20 1 r1_0_
rlabel metal3 569 10 569 10 1 r2_0_
rlabel metal3 571 120 571 120 1 r2_1_
rlabel metal3 571 130 571 130 1 r1_1
rlabel metal3 571 230 571 230 1 r2_2_
rlabel metal3 571 240 571 240 1 r1_2_
rlabel metal3 571 340 571 340 1 r2_3_
rlabel metal3 571 350 571 350 1 r1_3_
rlabel metal3 571 450 571 450 1 r2_4_
rlabel metal3 571 460 571 460 1 r1_4_
rlabel metal3 571 560 571 560 1 r2_5_
rlabel metal3 571 570 571 570 1 r1_5_
rlabel metal3 571 670 571 670 1 r2_6_
rlabel metal3 571 680 571 680 1 r1_6_
rlabel metal3 571 780 571 780 1 r2_7_
rlabel metal3 571 790 571 790 1 r1_7_
<< end >>
