magic
tech scmos
timestamp 1493149968
<< metal2 >>
rect 1135 1460 1138 1518
rect 1167 1470 1170 1519
rect 1199 1480 1202 1519
rect 1231 1490 1234 1517
rect 1295 1500 1298 1518
rect 1335 1510 1338 1519
rect 1321 1344 1325 1456
rect 1353 1342 1357 1466
rect 1529 1340 1533 1476
rect 1681 1344 1685 1486
rect 1713 1344 1717 1496
rect 1769 1344 1773 1506
rect 1937 1343 1941 1516
<< m3contact >>
rect 1366 1516 1370 1520
rect 1937 1516 1941 1520
rect 1335 1506 1339 1510
rect 1769 1506 1773 1510
rect 1295 1496 1299 1500
rect 1713 1496 1717 1500
rect 1231 1486 1235 1490
rect 1681 1486 1685 1490
rect 1199 1476 1203 1480
rect 1529 1476 1533 1480
rect 1167 1466 1171 1470
rect 1353 1466 1357 1470
rect 1135 1456 1139 1460
rect 1321 1456 1325 1460
<< metal3 >>
rect 1365 1520 1942 1521
rect 1365 1516 1366 1520
rect 1370 1516 1937 1520
rect 1941 1516 1942 1520
rect 1365 1515 1942 1516
rect 1334 1510 1774 1511
rect 1334 1506 1335 1510
rect 1339 1506 1769 1510
rect 1773 1506 1774 1510
rect 1334 1505 1774 1506
rect 1294 1500 1718 1501
rect 1294 1496 1295 1500
rect 1299 1496 1713 1500
rect 1717 1496 1718 1500
rect 1294 1495 1718 1496
rect 1230 1490 1686 1491
rect 1230 1486 1231 1490
rect 1235 1486 1681 1490
rect 1685 1486 1686 1490
rect 1230 1485 1686 1486
rect 1198 1480 1534 1481
rect 1198 1476 1199 1480
rect 1203 1476 1529 1480
rect 1533 1476 1534 1480
rect 1198 1475 1534 1476
rect 1166 1470 1358 1471
rect 1166 1466 1167 1470
rect 1171 1466 1353 1470
rect 1357 1466 1358 1470
rect 1166 1465 1358 1466
rect 1134 1460 1326 1461
rect 1134 1456 1135 1460
rect 1139 1456 1321 1460
rect 1325 1456 1326 1460
rect 1134 1455 1326 1456
use mips_fsm  mips_fsm_0
timestamp 1493147875
transform 1 0 965 0 1 1517
box 0 0 584 980
use datapath_new  datapath_new_0
timestamp 1493145788
transform 1 0 -279 0 1 32
box 279 -32 3123 2811
<< end >>
