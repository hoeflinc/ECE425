magic
tech scmos
timestamp 1492485052
<< metal1 >>
rect -47 1630 -1 1638
rect -47 1540 -1 1548
rect -26 1477 -8 1481
rect -26 1367 -15 1371
rect -41 1300 8 1308
rect -26 1257 -22 1261
rect -44 1210 5 1218
rect -45 1190 4 1198
rect -44 1100 5 1108
rect -41 1080 95 1088
rect -4 1040 1 1044
rect -40 970 96 978
rect -11 930 0 934
rect -41 860 95 868
rect -18 820 0 824
rect -41 770 95 778
rect -40 750 96 758
rect -25 710 0 714
rect -40 660 96 668
rect -40 640 96 648
rect -40 550 96 558
rect -41 530 95 538
rect -4 490 0 494
rect -42 440 94 448
rect -47 420 89 428
rect -11 380 0 384
rect -44 330 92 338
rect -43 310 93 318
rect -18 270 1 274
rect -43 220 93 228
rect -45 200 91 208
rect -25 160 1 164
rect -42 110 94 118
rect -44 90 92 98
rect -49 0 87 8
<< m2contact >>
rect -10 1644 -6 1648
rect 47 1644 51 1648
rect -28 1582 -24 1586
rect -8 1477 -4 1481
rect -15 1367 -11 1371
rect -22 1257 -18 1261
rect -29 1147 -25 1151
rect -1 1150 3 1154
rect -8 1040 -4 1044
rect -47 1030 -43 1034
rect -15 930 -11 934
rect -47 920 -43 924
rect -22 820 -18 824
rect -47 810 -43 814
rect 165 812 169 816
rect -29 710 -25 714
rect 165 702 169 706
rect -1 600 3 604
rect 165 592 169 596
rect -8 490 -4 494
rect 165 482 169 486
rect -15 380 -11 384
rect 165 372 169 376
rect -22 270 -18 274
rect 165 262 169 266
rect -29 160 -25 164
rect 165 152 169 156
rect -1 50 3 54
rect 165 42 169 46
<< metal2 >>
rect -28 1519 -24 1582
rect -2 1528 2 1563
rect -29 1145 -25 1147
rect -29 714 -25 1141
rect -22 824 -18 1257
rect -15 934 -11 1367
rect -8 1044 -4 1477
rect -1 1154 3 1515
rect 14 1324 18 1524
rect 14 1252 18 1320
rect 46 1246 50 1318
rect 14 1207 18 1239
rect 70 1208 74 1240
rect 78 1112 82 1320
rect 78 1032 82 1108
rect 126 1112 130 1113
rect -29 164 -25 591
rect -22 274 -18 701
rect -15 384 -11 811
rect -8 494 -4 921
rect -1 604 3 1031
rect 110 1026 114 1100
rect 78 988 82 1018
rect 126 922 130 1108
rect 134 988 138 1018
rect 158 916 162 992
rect 126 878 130 909
rect 182 878 186 913
rect -1 54 3 481
<< m3contact >>
rect -2 1524 2 1528
rect 14 1524 18 1528
rect -28 1515 -24 1519
rect -1 1515 3 1519
rect -29 1141 -25 1145
rect -47 1030 -43 1034
rect -47 920 -43 924
rect -171 812 -167 816
rect -47 810 -43 814
rect -164 725 -160 729
rect 14 1320 18 1324
rect 78 1320 82 1324
rect 14 1239 18 1243
rect 30 1239 34 1243
rect 30 1204 34 1208
rect 70 1204 74 1208
rect 78 1108 82 1112
rect -1 1031 3 1035
rect 126 1108 130 1112
rect -8 921 -4 925
rect -15 811 -11 815
rect -22 701 -18 705
rect -157 615 -153 619
rect -29 591 -25 595
rect -150 505 -146 509
rect -143 395 -139 399
rect -136 285 -132 289
rect -129 175 -125 179
rect 78 1018 82 1022
rect 94 1018 98 1022
rect 94 984 98 988
rect 134 984 138 988
rect 126 909 130 913
rect 142 909 146 913
rect 142 874 146 878
rect 182 874 186 878
rect -1 481 3 485
rect -122 65 -118 69
<< metal3 >>
rect -3 1528 19 1529
rect -3 1524 -2 1528
rect 2 1524 14 1528
rect 18 1524 19 1528
rect -3 1523 19 1524
rect -29 1519 4 1520
rect -29 1515 -28 1519
rect -24 1515 -1 1519
rect 3 1515 4 1519
rect -29 1514 4 1515
rect 13 1324 83 1325
rect 13 1320 14 1324
rect 18 1320 78 1324
rect 82 1320 83 1324
rect 13 1319 83 1320
rect 13 1243 35 1244
rect 13 1239 14 1243
rect 18 1239 30 1243
rect 34 1239 35 1243
rect 13 1238 35 1239
rect 29 1208 75 1209
rect 29 1204 30 1208
rect 34 1204 70 1208
rect 74 1204 75 1208
rect 29 1203 75 1204
rect -30 1145 1 1146
rect -30 1141 -29 1145
rect -25 1141 1 1145
rect -30 1140 1 1141
rect 77 1112 131 1113
rect 77 1108 78 1112
rect 82 1108 126 1112
rect 130 1108 131 1112
rect 77 1107 131 1108
rect -48 1035 0 1036
rect -48 1034 -1 1035
rect -48 1030 -47 1034
rect -43 1031 -1 1034
rect -43 1030 0 1031
rect -48 1029 0 1030
rect 77 1022 99 1023
rect 77 1018 78 1022
rect 82 1018 94 1022
rect 98 1018 99 1022
rect 77 1017 99 1018
rect 93 988 139 989
rect 93 984 94 988
rect 98 984 134 988
rect 138 984 139 988
rect 93 983 139 984
rect -48 925 0 926
rect -48 924 -8 925
rect -48 920 -47 924
rect -43 921 -8 924
rect -4 921 0 925
rect -43 920 0 921
rect -48 919 0 920
rect 125 913 147 914
rect 125 909 126 913
rect 130 909 142 913
rect 146 909 147 913
rect 125 908 147 909
rect 141 878 187 879
rect 141 874 142 878
rect 146 874 182 878
rect 186 874 187 878
rect 141 873 187 874
rect -48 815 0 816
rect -48 814 -15 815
rect -48 810 -47 814
rect -43 811 -15 814
rect -11 811 0 815
rect -43 810 0 811
rect -48 809 0 810
rect -28 705 1 706
rect -28 701 -22 705
rect -18 701 1 705
rect -28 700 1 701
rect -27 595 2 596
rect -25 591 2 595
rect -27 590 2 591
rect -28 485 1 486
rect -28 481 -1 485
rect -28 480 1 481
rect -28 370 1 376
rect -29 260 0 266
rect -28 150 1 156
rect -28 40 1 46
use xor2_2x  xor2_2x_0
timestamp 1492457336
transform 1 0 6 0 1 1214
box -6 -4 74 96
use xor2_2x  xor2_2x_1
timestamp 1492457336
transform 1 0 70 0 1 994
box -6 -4 74 96
use shift_source_gen  shift_source_gen_0
timestamp 1492473219
transform 1 0 -74 0 1 0
box -98 0 162 1648
use xor2_2x  xor2_2x_2
timestamp 1492457336
transform 1 0 118 0 1 884
box -6 -4 74 96
use log_shifter  log_shifter_0
timestamp 1492474365
transform 1 0 112 0 1 0
box -112 0 57 1208
<< labels >>
rlabel metal2 48 1316 48 1316 1 s2
rlabel metal2 112 1098 112 1098 1 s1
rlabel metal2 160 990 160 990 1 s0
rlabel m2contact -8 1648 -8 1648 5 right
rlabel m3contact -120 67 -120 67 1 a0
rlabel m3contact -127 177 -127 177 1 a1
rlabel m3contact -134 287 -134 287 1 a2
rlabel m3contact -141 397 -141 397 1 a3
rlabel m3contact -148 507 -148 507 1 a4
rlabel m3contact -155 617 -155 617 1 a5
rlabel m3contact -162 727 -162 727 1 a6
rlabel m3contact -169 814 -169 814 3 a7
rlabel m2contact 167 704 167 704 1 y6
rlabel m2contact 167 814 167 814 1 y7
rlabel m2contact 167 594 167 594 1 y5
rlabel m2contact 167 484 167 484 1 y4
rlabel m2contact 167 374 167 374 1 y3
rlabel m2contact 167 264 167 264 1 y2
rlabel m2contact 167 154 167 154 1 y1
rlabel m2contact 167 44 167 44 1 y0
rlabel m2contact 49 1646 49 1646 5 arith
rlabel m2contact 49 1648 49 1648 5 arith
rlabel metal3 -16 44 -16 44 1 z0
rlabel metal3 -15 154 -15 154 1 z1
rlabel metal3 144 873 144 873 1 s0xor
rlabel metal3 -14 263 -14 263 1 z2
rlabel metal3 -13 373 -13 373 1 z3
rlabel metal3 -14 483 -14 483 1 z4
rlabel metal3 -9 594 -9 594 1 z5
rlabel metal3 -9 704 -9 704 1 z6
rlabel metal3 -21 812 -21 812 1 z7
rlabel metal3 -11 923 -11 923 1 z8
rlabel metal3 -4 1032 -4 1032 1 z9
rlabel metal3 -24 1143 -24 1143 1 z10
rlabel metal1 -24 1259 -24 1259 1 z11
rlabel metal1 -19 1368 -19 1368 1 z12
rlabel metal1 -18 1479 -18 1479 1 z13
rlabel metal2 -25 1575 -25 1575 1 z14
<< end >>
