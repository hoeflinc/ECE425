magic
tech scmos
timestamp 1492465660
<< metal1 >>
rect 31 1582 46 1586
<< m2contact >>
rect 46 1582 50 1586
<< metal2 >>
rect -41 1476 -37 1582
rect -41 1366 -37 1472
rect -41 1256 -37 1362
rect -69 509 -65 1155
rect -41 1146 -37 1252
rect -62 289 -58 1045
rect -41 1036 -37 1142
rect -55 179 -51 935
rect -41 926 -37 1032
rect -48 69 -44 825
rect -41 816 -37 922
rect -34 1563 -30 1583
rect -34 809 -30 1559
rect -10 1553 -6 1583
rect -2 1567 2 1594
rect 14 1567 18 1603
rect 64 1582 68 1648
rect 121 1605 125 1648
rect 72 1567 76 1586
rect 88 1565 92 1586
rect 14 1556 18 1561
rect 112 1565 116 1578
rect -10 919 -6 1549
rect 88 1537 92 1561
rect 152 1553 156 1586
rect -10 767 -6 813
rect 38 767 42 1533
rect -10 763 42 767
rect 22 34 26 763
<< m3contact >>
rect -41 1582 -37 1586
rect -41 1472 -37 1476
rect -41 1362 -37 1366
rect -41 1252 -37 1256
rect -69 1155 -65 1159
rect -41 1142 -37 1146
rect -69 505 -65 509
rect -62 1045 -58 1049
rect -41 1032 -37 1036
rect -62 285 -58 289
rect -55 935 -51 939
rect -41 922 -37 926
rect -55 175 -51 179
rect -48 825 -44 829
rect -41 812 -37 816
rect -34 1559 -30 1563
rect 96 1582 100 1586
rect 128 1582 132 1586
rect 72 1559 76 1563
rect 88 1561 92 1565
rect 112 1561 116 1565
rect -10 1549 -6 1553
rect 152 1549 156 1553
rect 38 1533 42 1537
rect 88 1533 92 1537
rect -48 65 -44 69
rect 31 725 35 729
rect 31 615 35 619
rect 31 505 35 509
rect 31 395 35 399
rect 31 285 35 289
rect 31 175 35 179
rect 31 65 35 69
<< metal3 >>
rect 95 1586 133 1587
rect 95 1582 96 1586
rect 100 1582 128 1586
rect 132 1582 133 1586
rect 95 1581 133 1582
rect 87 1565 117 1566
rect -35 1563 77 1564
rect -35 1559 -34 1563
rect -30 1559 72 1563
rect 76 1559 77 1563
rect 87 1561 88 1565
rect 92 1561 112 1565
rect 116 1561 117 1565
rect 87 1560 117 1561
rect -35 1558 77 1559
rect -11 1553 157 1554
rect -11 1549 -10 1553
rect -6 1549 152 1553
rect 156 1549 157 1553
rect -11 1548 157 1549
rect 37 1537 93 1538
rect 37 1533 38 1537
rect 42 1533 88 1537
rect 92 1533 93 1537
rect 37 1532 93 1533
rect -70 1159 -49 1160
rect -70 1155 -69 1159
rect -65 1155 -49 1159
rect -70 1154 -49 1155
rect -63 1049 -49 1050
rect -63 1045 -62 1049
rect -58 1045 -49 1049
rect -63 1044 -49 1045
rect -56 939 -49 940
rect -56 935 -55 939
rect -51 935 -49 939
rect -56 934 -49 935
rect -13 729 36 730
rect -13 725 31 729
rect 35 725 36 729
rect -13 724 36 725
rect -13 619 36 620
rect -13 615 31 619
rect 35 615 36 619
rect -13 614 36 615
rect -70 509 36 510
rect -70 505 -69 509
rect -65 505 31 509
rect 35 505 36 509
rect -70 504 36 505
rect -13 399 36 400
rect -13 395 31 399
rect 35 395 36 399
rect -13 394 36 395
rect -63 289 36 290
rect -63 285 -62 289
rect -58 285 31 289
rect 35 285 36 289
rect -63 284 36 285
rect -56 179 36 180
rect -56 175 -55 179
rect -51 175 31 179
rect 35 175 36 179
rect -56 174 36 175
rect -49 69 36 70
rect -49 65 -48 69
rect -44 65 31 69
rect 35 65 36 69
rect -49 64 36 65
use nandnandnand_1x  nandnandnand_1x_0
array 1 1 80 1 8 110
timestamp 1492464959
transform 1 0 -40 0 1 770
box -9 0 80 100
use invbuf_4x  invbuf_4x_1
timestamp 1484532969
transform 1 0 64 0 1 1544
box -6 -4 34 96
use and2_1x  and2_1x_1
timestamp 1484419738
transform 1 0 96 0 1 1544
box -6 -4 34 96
use invbuf_4x  invbuf_4x_0
timestamp 1484532969
transform 1 0 128 0 1 1544
box -6 -4 34 96
use and2_1x  and2_1x_0
array 0 0 40 1 7 110
timestamp 1484419738
transform 1 0 6 0 1 4
box -6 -4 34 96
<< labels >>
rlabel metal2 66 1646 66 1646 5 right
rlabel metal2 123 1646 123 1646 5 arith
<< end >>
