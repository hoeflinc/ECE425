magic
tech scmos
timestamp 1488306862
<< m2contact >>
rect -7 -2 7 2
<< end >>
