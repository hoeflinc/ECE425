magic
tech scmos
timestamp 1493745683
<< m2contact >>
rect -7 -7 7 7
<< end >>
