magic
tech scmos
timestamp 1493745683
<< m2contact >>
rect -2 -2 2 2
<< end >>
