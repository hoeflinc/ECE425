magic
tech scmos
timestamp 1486492580
<< nwell >>
rect -6 40 34 96
<< ntransistor >>
rect 5 6 7 22
rect 10 6 12 22
rect 15 6 17 22
<< ptransistor >>
rect 5 69 7 82
rect 13 69 15 82
rect 21 69 23 82
<< ndiffusion >>
rect 0 20 5 22
rect 4 8 5 20
rect 0 6 5 8
rect 7 6 10 22
rect 12 6 15 22
rect 17 20 22 22
rect 17 8 18 20
rect 17 6 22 8
<< pdiffusion >>
rect 0 81 5 82
rect 4 69 5 81
rect 7 81 13 82
rect 7 69 8 81
rect 12 69 13 81
rect 15 81 21 82
rect 15 69 16 81
rect 20 69 21 81
rect 23 81 28 82
rect 23 69 24 81
<< ndcontact >>
rect 0 8 4 20
rect 18 8 22 20
<< pdcontact >>
rect 0 69 4 81
rect 8 69 12 81
rect 16 69 20 81
rect 24 69 28 81
<< psubstratepcontact >>
rect 0 -2 4 2
rect 8 -2 12 2
rect 16 -2 20 2
rect 24 -2 28 2
<< nsubstratencontact >>
rect 0 88 4 92
rect 8 88 12 92
rect 16 88 20 92
rect 24 88 28 92
<< polysilicon >>
rect 5 82 7 84
rect 13 82 15 84
rect 21 82 23 84
rect 5 65 7 69
rect 13 65 15 69
rect 1 63 7 65
rect 10 63 15 65
rect 1 47 3 63
rect 10 47 12 63
rect 21 58 23 69
rect 20 56 23 58
rect 1 25 3 43
rect 1 23 7 25
rect 5 22 7 23
rect 10 22 12 43
rect 20 25 22 56
rect 15 23 22 25
rect 15 22 17 23
rect 5 4 7 6
rect 10 4 12 6
rect 15 4 17 6
<< polycontact >>
rect 0 43 4 47
rect 8 43 12 47
rect 16 43 20 47
<< metal1 >>
rect -2 92 30 94
rect -2 88 0 92
rect 4 88 8 92
rect 12 88 16 92
rect 20 88 24 92
rect 28 88 30 92
rect -2 86 30 88
rect 0 81 4 86
rect 16 81 20 86
rect 8 63 12 69
rect 24 63 28 69
rect 8 59 28 63
rect 24 47 28 59
rect 24 21 28 43
rect 0 20 4 21
rect 22 17 28 21
rect 0 4 4 8
rect -2 2 30 4
rect -2 -2 0 2
rect 4 -2 8 2
rect 12 -2 16 2
rect 20 -2 24 2
rect 28 -2 30 2
rect -2 -4 30 -2
<< m2contact >>
rect 0 43 4 47
rect 8 43 12 47
rect 16 43 20 47
rect 24 43 28 47
<< labels >>
rlabel metal1 0 0 0 0 1 Gnd!
rlabel metal1 -1 90 -1 90 3 Vdd!
rlabel m2contact 10 45 10 45 1 B
rlabel m2contact 18 45 18 45 1 C
rlabel m2contact 26 45 26 45 1 Y
rlabel m2contact 2 45 2 45 1 A
<< end >>
